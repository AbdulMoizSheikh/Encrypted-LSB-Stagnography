magic
tech sky130A
magscale 1 2
timestamp 1661348181
<< checkpaint >>
rect -12658 -11586 596582 715522
<< locali >>
rect 239229 456943 239263 457249
rect 255053 457011 255087 457249
rect 266093 457147 266127 457249
rect 283481 456875 283515 457453
rect 377597 456807 377631 457385
rect 379161 457215 379195 457385
rect 380909 457079 380943 457385
rect 288265 336447 288299 336549
rect 283205 335971 283239 336277
rect 293417 335631 293451 336413
rect 354597 336243 354631 336413
rect 378701 335767 378735 336413
rect 378793 335903 378827 336481
rect 382289 336243 382323 336549
rect 393237 336107 393271 336413
rect 393179 336073 393271 336107
rect 413109 335359 413143 335597
rect 414799 335597 415225 335631
rect 414489 335359 414523 335597
rect 414581 335359 414615 335529
rect 387165 335223 387199 335325
rect 407865 333183 407899 333353
rect 258123 8109 258457 8143
rect 258089 7871 258123 7973
rect 53941 3383 53975 3621
rect 84393 3383 84427 4029
rect 317889 3961 318199 3995
rect 317889 3587 317923 3961
rect 318165 3927 318199 3961
rect 318073 3791 318107 3893
rect 317981 3587 318015 3757
rect 320373 3519 320407 3893
rect 358645 3825 358921 3859
rect 358645 3791 358679 3825
rect 329021 3587 329055 3757
rect 329205 3451 329239 3553
rect 535009 3383 535043 4097
rect 102149 3179 102183 3281
rect 102091 3145 102183 3179
rect 111165 2907 111199 3077
rect 354229 3043 354263 3145
rect 122205 2771 122239 2873
rect 125551 2805 125701 2839
rect 122205 2737 122389 2771
<< viali >>
rect 283481 457453 283515 457487
rect 239229 457249 239263 457283
rect 255053 457249 255087 457283
rect 266093 457249 266127 457283
rect 266093 457113 266127 457147
rect 255053 456977 255087 457011
rect 239229 456909 239263 456943
rect 283481 456841 283515 456875
rect 377597 457385 377631 457419
rect 379161 457385 379195 457419
rect 379161 457181 379195 457215
rect 380909 457385 380943 457419
rect 380909 457045 380943 457079
rect 377597 456773 377631 456807
rect 288265 336549 288299 336583
rect 382289 336549 382323 336583
rect 378793 336481 378827 336515
rect 288265 336413 288299 336447
rect 293417 336413 293451 336447
rect 283205 336277 283239 336311
rect 283205 335937 283239 335971
rect 354597 336413 354631 336447
rect 354597 336209 354631 336243
rect 378701 336413 378735 336447
rect 382289 336209 382323 336243
rect 393237 336413 393271 336447
rect 393145 336073 393179 336107
rect 378793 335869 378827 335903
rect 378701 335733 378735 335767
rect 293417 335597 293451 335631
rect 413109 335597 413143 335631
rect 387165 335325 387199 335359
rect 413109 335325 413143 335359
rect 414489 335597 414523 335631
rect 414765 335597 414799 335631
rect 415225 335597 415259 335631
rect 414489 335325 414523 335359
rect 414581 335529 414615 335563
rect 414581 335325 414615 335359
rect 387165 335189 387199 335223
rect 407865 333353 407899 333387
rect 407865 333149 407899 333183
rect 258089 8109 258123 8143
rect 258457 8109 258491 8143
rect 258089 7973 258123 8007
rect 258089 7837 258123 7871
rect 535009 4097 535043 4131
rect 84393 4029 84427 4063
rect 53941 3621 53975 3655
rect 53941 3349 53975 3383
rect 318073 3893 318107 3927
rect 318165 3893 318199 3927
rect 320373 3893 320407 3927
rect 317889 3553 317923 3587
rect 317981 3757 318015 3791
rect 318073 3757 318107 3791
rect 317981 3553 318015 3587
rect 358921 3825 358955 3859
rect 329021 3757 329055 3791
rect 358645 3757 358679 3791
rect 329021 3553 329055 3587
rect 329205 3553 329239 3587
rect 320373 3485 320407 3519
rect 329205 3417 329239 3451
rect 84393 3349 84427 3383
rect 535009 3349 535043 3383
rect 102149 3281 102183 3315
rect 102057 3145 102091 3179
rect 354229 3145 354263 3179
rect 111165 3077 111199 3111
rect 354229 3009 354263 3043
rect 111165 2873 111199 2907
rect 122205 2873 122239 2907
rect 125517 2805 125551 2839
rect 125701 2805 125735 2839
rect 122389 2737 122423 2771
<< metal1 >>
rect 317322 700952 317328 701004
rect 317380 700992 317386 701004
rect 429838 700992 429844 701004
rect 317380 700964 429844 700992
rect 317380 700952 317386 700964
rect 429838 700952 429844 700964
rect 429896 700952 429902 701004
rect 202782 700884 202788 700936
rect 202840 700924 202846 700936
rect 331306 700924 331312 700936
rect 202840 700896 331312 700924
rect 202840 700884 202846 700896
rect 331306 700884 331312 700896
rect 331364 700884 331370 700936
rect 313182 700816 313188 700868
rect 313240 700856 313246 700868
rect 462314 700856 462320 700868
rect 313240 700828 462320 700856
rect 313240 700816 313246 700828
rect 462314 700816 462320 700828
rect 462372 700816 462378 700868
rect 315942 700748 315948 700800
rect 316000 700788 316006 700800
rect 478506 700788 478512 700800
rect 316000 700760 478512 700788
rect 316000 700748 316006 700760
rect 478506 700748 478512 700760
rect 478564 700748 478570 700800
rect 311802 700680 311808 700732
rect 311860 700720 311866 700732
rect 494790 700720 494796 700732
rect 311860 700692 494796 700720
rect 311860 700680 311866 700692
rect 494790 700680 494796 700692
rect 494848 700680 494854 700732
rect 137830 700612 137836 700664
rect 137888 700652 137894 700664
rect 336734 700652 336740 700664
rect 137888 700624 336740 700652
rect 137888 700612 137894 700624
rect 336734 700612 336740 700624
rect 336792 700612 336798 700664
rect 309042 700544 309048 700596
rect 309100 700584 309106 700596
rect 527174 700584 527180 700596
rect 309100 700556 527180 700584
rect 309100 700544 309106 700556
rect 527174 700544 527180 700556
rect 527232 700544 527238 700596
rect 105446 700476 105452 700528
rect 105504 700516 105510 700528
rect 106182 700516 106188 700528
rect 105504 700488 106188 700516
rect 105504 700476 105510 700488
rect 106182 700476 106188 700488
rect 106240 700476 106246 700528
rect 310422 700476 310428 700528
rect 310480 700516 310486 700528
rect 543458 700516 543464 700528
rect 310480 700488 543464 700516
rect 310480 700476 310486 700488
rect 543458 700476 543464 700488
rect 543516 700476 543522 700528
rect 40494 700408 40500 700460
rect 40552 700448 40558 700460
rect 41322 700448 41328 700460
rect 40552 700420 41328 700448
rect 40552 700408 40558 700420
rect 41322 700408 41328 700420
rect 41380 700408 41386 700460
rect 307662 700408 307668 700460
rect 307720 700448 307726 700460
rect 559650 700448 559656 700460
rect 307720 700420 559656 700448
rect 307720 700408 307726 700420
rect 559650 700408 559656 700420
rect 559708 700408 559714 700460
rect 72970 700340 72976 700392
rect 73028 700380 73034 700392
rect 340874 700380 340880 700392
rect 73028 700352 340880 700380
rect 73028 700340 73034 700352
rect 340874 700340 340880 700352
rect 340932 700340 340938 700392
rect 8110 700272 8116 700324
rect 8168 700312 8174 700324
rect 345014 700312 345020 700324
rect 8168 700284 345020 700312
rect 8168 700272 8174 700284
rect 345014 700272 345020 700284
rect 345072 700272 345078 700324
rect 320082 700204 320088 700256
rect 320140 700244 320146 700256
rect 413646 700244 413652 700256
rect 320140 700216 413652 700244
rect 320140 700204 320146 700216
rect 413646 700204 413652 700216
rect 413704 700204 413710 700256
rect 318702 700136 318708 700188
rect 318760 700176 318766 700188
rect 397454 700176 397460 700188
rect 318760 700148 397460 700176
rect 318760 700136 318766 700148
rect 397454 700136 397460 700148
rect 397512 700136 397518 700188
rect 267642 700068 267648 700120
rect 267700 700108 267706 700120
rect 327074 700108 327080 700120
rect 267700 700080 327080 700108
rect 267700 700068 267706 700080
rect 327074 700068 327080 700080
rect 327132 700068 327138 700120
rect 321462 700000 321468 700052
rect 321520 700040 321526 700052
rect 364978 700040 364984 700052
rect 321520 700012 364984 700040
rect 321520 700000 321526 700012
rect 364978 700000 364984 700012
rect 365036 700000 365042 700052
rect 324222 699932 324228 699984
rect 324280 699972 324286 699984
rect 348786 699972 348792 699984
rect 324280 699944 348792 699972
rect 324280 699932 324286 699944
rect 348786 699932 348792 699944
rect 348844 699932 348850 699984
rect 322842 699864 322848 699916
rect 322900 699904 322906 699916
rect 332502 699904 332508 699916
rect 322900 699876 332508 699904
rect 322900 699864 322906 699876
rect 332502 699864 332508 699876
rect 332560 699864 332566 699916
rect 24302 699660 24308 699712
rect 24360 699700 24366 699712
rect 24762 699700 24768 699712
rect 24360 699672 24768 699700
rect 24360 699660 24366 699672
rect 24762 699660 24768 699672
rect 24820 699660 24826 699712
rect 170306 699660 170312 699712
rect 170364 699700 170370 699712
rect 171042 699700 171048 699712
rect 170364 699672 171048 699700
rect 170364 699660 170370 699672
rect 171042 699660 171048 699672
rect 171100 699660 171106 699712
rect 235166 699660 235172 699712
rect 235224 699700 235230 699712
rect 235902 699700 235908 699712
rect 235224 699672 235908 699700
rect 235224 699660 235230 699672
rect 235902 699660 235908 699672
rect 235960 699660 235966 699712
rect 300118 699660 300124 699712
rect 300176 699700 300182 699712
rect 300762 699700 300768 699712
rect 300176 699672 300768 699700
rect 300176 699660 300182 699672
rect 300762 699660 300768 699672
rect 300820 699660 300826 699712
rect 304902 696940 304908 696992
rect 304960 696980 304966 696992
rect 580166 696980 580172 696992
rect 304960 696952 580172 696980
rect 304960 696940 304966 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 306282 683136 306288 683188
rect 306340 683176 306346 683188
rect 580166 683176 580172 683188
rect 306340 683148 580172 683176
rect 306340 683136 306346 683148
rect 580166 683136 580172 683148
rect 580224 683136 580230 683188
rect 302142 670760 302148 670812
rect 302200 670800 302206 670812
rect 580166 670800 580172 670812
rect 302200 670772 580172 670800
rect 302200 670760 302206 670772
rect 580166 670760 580172 670772
rect 580224 670760 580230 670812
rect 3510 670692 3516 670744
rect 3568 670732 3574 670744
rect 333238 670732 333244 670744
rect 3568 670704 333244 670732
rect 3568 670692 3574 670704
rect 333238 670692 333244 670704
rect 333296 670692 333302 670744
rect 3510 656888 3516 656940
rect 3568 656928 3574 656940
rect 350534 656928 350540 656940
rect 3568 656900 350540 656928
rect 3568 656888 3574 656900
rect 350534 656888 350540 656900
rect 350592 656888 350598 656940
rect 299382 643084 299388 643136
rect 299440 643124 299446 643136
rect 580166 643124 580172 643136
rect 299440 643096 580172 643124
rect 299440 643084 299446 643096
rect 580166 643084 580172 643096
rect 580224 643084 580230 643136
rect 300670 630640 300676 630692
rect 300728 630680 300734 630692
rect 580166 630680 580172 630692
rect 300728 630652 580172 630680
rect 300728 630640 300734 630652
rect 580166 630640 580172 630652
rect 580224 630640 580230 630692
rect 3326 618264 3332 618316
rect 3384 618304 3390 618316
rect 338758 618304 338764 618316
rect 3384 618276 338764 618304
rect 3384 618264 3390 618276
rect 338758 618264 338764 618276
rect 338816 618264 338822 618316
rect 298002 616836 298008 616888
rect 298060 616876 298066 616888
rect 580166 616876 580172 616888
rect 298060 616848 580172 616876
rect 298060 616836 298066 616848
rect 580166 616836 580172 616848
rect 580224 616836 580230 616888
rect 3326 605820 3332 605872
rect 3384 605860 3390 605872
rect 354674 605860 354680 605872
rect 3384 605832 354680 605860
rect 3384 605820 3390 605832
rect 354674 605820 354680 605832
rect 354732 605820 354738 605872
rect 295242 590656 295248 590708
rect 295300 590696 295306 590708
rect 579798 590696 579804 590708
rect 295300 590668 579804 590696
rect 295300 590656 295306 590668
rect 579798 590656 579804 590668
rect 579856 590656 579862 590708
rect 296622 576852 296628 576904
rect 296680 576892 296686 576904
rect 580166 576892 580172 576904
rect 296680 576864 580172 576892
rect 296680 576852 296686 576864
rect 580166 576852 580172 576864
rect 580224 576852 580230 576904
rect 3050 565836 3056 565888
rect 3108 565876 3114 565888
rect 342898 565876 342904 565888
rect 3108 565848 342904 565876
rect 3108 565836 3114 565848
rect 342898 565836 342904 565848
rect 342956 565836 342962 565888
rect 293862 563048 293868 563100
rect 293920 563088 293926 563100
rect 579798 563088 579804 563100
rect 293920 563060 579804 563088
rect 293920 563048 293926 563060
rect 579798 563048 579804 563060
rect 579856 563048 579862 563100
rect 3326 553392 3332 553444
rect 3384 553432 3390 553444
rect 360194 553432 360200 553444
rect 3384 553404 360200 553432
rect 3384 553392 3390 553404
rect 360194 553392 360200 553404
rect 360252 553392 360258 553444
rect 289722 536800 289728 536852
rect 289780 536840 289786 536852
rect 580166 536840 580172 536852
rect 289780 536812 580172 536840
rect 289780 536800 289786 536812
rect 580166 536800 580172 536812
rect 580224 536800 580230 536852
rect 291102 524424 291108 524476
rect 291160 524464 291166 524476
rect 580166 524464 580172 524476
rect 291160 524436 580172 524464
rect 291160 524424 291166 524436
rect 580166 524424 580172 524436
rect 580224 524424 580230 524476
rect 3326 514768 3332 514820
rect 3384 514808 3390 514820
rect 348418 514808 348424 514820
rect 3384 514780 348424 514808
rect 3384 514768 3390 514780
rect 348418 514768 348424 514780
rect 348476 514768 348482 514820
rect 288342 510620 288348 510672
rect 288400 510660 288406 510672
rect 580166 510660 580172 510672
rect 288400 510632 580172 510660
rect 288400 510620 288406 510632
rect 580166 510620 580172 510632
rect 580224 510620 580230 510672
rect 3234 500964 3240 501016
rect 3292 501004 3298 501016
rect 364334 501004 364340 501016
rect 3292 500976 364340 501004
rect 3292 500964 3298 500976
rect 364334 500964 364340 500976
rect 364392 500964 364398 501016
rect 285582 484372 285588 484424
rect 285640 484412 285646 484424
rect 580166 484412 580172 484424
rect 285640 484384 580172 484412
rect 285640 484372 285646 484384
rect 580166 484372 580172 484384
rect 580224 484372 580230 484424
rect 286962 470568 286968 470620
rect 287020 470608 287026 470620
rect 579982 470608 579988 470620
rect 287020 470580 579988 470608
rect 287020 470568 287026 470580
rect 579982 470568 579988 470580
rect 580040 470568 580046 470620
rect 3510 462340 3516 462392
rect 3568 462380 3574 462392
rect 352558 462380 352564 462392
rect 3568 462352 352564 462380
rect 3568 462340 3574 462352
rect 352558 462340 352564 462352
rect 352616 462340 352622 462392
rect 171042 460844 171048 460896
rect 171100 460884 171106 460896
rect 334894 460884 334900 460896
rect 171100 460856 334900 460884
rect 171100 460844 171106 460856
rect 334894 460844 334900 460856
rect 334952 460844 334958 460896
rect 154482 460776 154488 460828
rect 154540 460816 154546 460828
rect 338114 460816 338120 460828
rect 154540 460788 338120 460816
rect 154540 460776 154546 460788
rect 338114 460776 338120 460788
rect 338172 460776 338178 460828
rect 338758 460776 338764 460828
rect 338816 460816 338822 460828
rect 356974 460816 356980 460828
rect 338816 460788 356980 460816
rect 338816 460776 338822 460788
rect 356974 460776 356980 460788
rect 357032 460776 357038 460828
rect 106182 460708 106188 460760
rect 106240 460748 106246 460760
rect 339678 460748 339684 460760
rect 106240 460720 339684 460748
rect 106240 460708 106246 460720
rect 339678 460708 339684 460720
rect 339736 460708 339742 460760
rect 89622 460640 89628 460692
rect 89680 460680 89686 460692
rect 342806 460680 342812 460692
rect 89680 460652 342812 460680
rect 89680 460640 89686 460652
rect 342806 460640 342812 460652
rect 342864 460640 342870 460692
rect 342898 460640 342904 460692
rect 342956 460680 342962 460692
rect 361758 460680 361764 460692
rect 342956 460652 361764 460680
rect 342956 460640 342962 460652
rect 361758 460640 361764 460652
rect 361816 460640 361822 460692
rect 41322 460572 41328 460624
rect 41380 460612 41386 460624
rect 344370 460612 344376 460624
rect 41380 460584 344376 460612
rect 41380 460572 41386 460584
rect 344370 460572 344376 460584
rect 344428 460572 344434 460624
rect 24762 460504 24768 460556
rect 24820 460544 24826 460556
rect 347774 460544 347780 460556
rect 24820 460516 347780 460544
rect 24820 460504 24826 460516
rect 347774 460504 347780 460516
rect 347832 460504 347838 460556
rect 348418 460504 348424 460556
rect 348476 460544 348482 460556
rect 366450 460544 366456 460556
rect 348476 460516 366456 460544
rect 348476 460504 348482 460516
rect 366450 460504 366456 460516
rect 366508 460504 366514 460556
rect 3418 460436 3424 460488
rect 3476 460476 3482 460488
rect 349154 460476 349160 460488
rect 3476 460448 349160 460476
rect 3476 460436 3482 460448
rect 349154 460436 349160 460448
rect 349212 460436 349218 460488
rect 352558 460436 352564 460488
rect 352616 460476 352622 460488
rect 371234 460476 371240 460488
rect 352616 460448 371240 460476
rect 352616 460436 352622 460448
rect 371234 460436 371240 460448
rect 371292 460436 371298 460488
rect 3602 460368 3608 460420
rect 3660 460408 3666 460420
rect 353846 460408 353852 460420
rect 3660 460380 353852 460408
rect 3660 460368 3666 460380
rect 353846 460368 353852 460380
rect 353904 460368 353910 460420
rect 3694 460300 3700 460352
rect 3752 460340 3758 460352
rect 358814 460340 358820 460352
rect 3752 460312 358820 460340
rect 3752 460300 3758 460312
rect 358814 460300 358820 460312
rect 358872 460300 358878 460352
rect 3786 460232 3792 460284
rect 3844 460272 3850 460284
rect 363322 460272 363328 460284
rect 3844 460244 363328 460272
rect 3844 460232 3850 460244
rect 363322 460232 363328 460244
rect 363380 460232 363386 460284
rect 3878 460164 3884 460216
rect 3936 460204 3942 460216
rect 368106 460204 368112 460216
rect 3936 460176 368112 460204
rect 3936 460164 3942 460176
rect 368106 460164 368112 460176
rect 368164 460164 368170 460216
rect 219342 460096 219348 460148
rect 219400 460136 219406 460148
rect 219400 460108 333192 460136
rect 219400 460096 219406 460108
rect 235902 460028 235908 460080
rect 235960 460068 235966 460080
rect 330202 460068 330208 460080
rect 235960 460040 330208 460068
rect 235960 460028 235966 460040
rect 330202 460028 330208 460040
rect 330260 460028 330266 460080
rect 333164 460068 333192 460108
rect 333238 460096 333244 460148
rect 333296 460136 333302 460148
rect 352282 460136 352288 460148
rect 333296 460108 352288 460136
rect 333296 460096 333302 460108
rect 352282 460096 352288 460108
rect 352340 460096 352346 460148
rect 333330 460068 333336 460080
rect 333164 460040 333336 460068
rect 333330 460028 333336 460040
rect 333388 460028 333394 460080
rect 284202 459960 284208 460012
rect 284260 460000 284266 460012
rect 328546 460000 328552 460012
rect 284260 459972 328552 460000
rect 284260 459960 284266 459972
rect 328546 459960 328552 459972
rect 328604 459960 328610 460012
rect 325694 459932 325700 459944
rect 316006 459904 325700 459932
rect 300762 459824 300768 459876
rect 300820 459864 300826 459876
rect 316006 459864 316034 459904
rect 325694 459892 325700 459904
rect 325752 459892 325758 459944
rect 300820 459836 316034 459864
rect 300820 459824 300826 459836
rect 281442 459756 281448 459808
rect 281500 459796 281506 459808
rect 281500 459768 287054 459796
rect 281500 459756 281506 459768
rect 285030 459688 285036 459740
rect 285088 459728 285094 459740
rect 285582 459728 285588 459740
rect 285088 459700 285588 459728
rect 285088 459688 285094 459700
rect 285582 459688 285588 459700
rect 285640 459688 285646 459740
rect 287026 459728 287054 459768
rect 292942 459756 292948 459808
rect 293000 459796 293006 459808
rect 293862 459796 293868 459808
rect 293000 459768 293868 459796
rect 293000 459756 293006 459768
rect 293862 459756 293868 459768
rect 293920 459756 293926 459808
rect 294506 459756 294512 459808
rect 294564 459796 294570 459808
rect 295242 459796 295248 459808
rect 294564 459768 295248 459796
rect 294564 459756 294570 459768
rect 295242 459756 295248 459768
rect 295300 459756 295306 459808
rect 296070 459756 296076 459808
rect 296128 459796 296134 459808
rect 296622 459796 296628 459808
rect 296128 459768 296628 459796
rect 296128 459756 296134 459768
rect 296622 459756 296628 459768
rect 296680 459756 296686 459808
rect 303982 459756 303988 459808
rect 304040 459796 304046 459808
rect 304902 459796 304908 459808
rect 304040 459768 304908 459796
rect 304040 459756 304046 459768
rect 304902 459756 304908 459768
rect 304960 459756 304966 459808
rect 305546 459756 305552 459808
rect 305604 459796 305610 459808
rect 306282 459796 306288 459808
rect 305604 459768 306288 459796
rect 305604 459756 305610 459768
rect 306282 459756 306288 459768
rect 306340 459756 306346 459808
rect 307110 459756 307116 459808
rect 307168 459796 307174 459808
rect 307662 459796 307668 459808
rect 307168 459768 307668 459796
rect 307168 459756 307174 459768
rect 307662 459756 307668 459768
rect 307720 459756 307726 459808
rect 315022 459756 315028 459808
rect 315080 459796 315086 459808
rect 315942 459796 315948 459808
rect 315080 459768 315948 459796
rect 315080 459756 315086 459768
rect 315942 459756 315948 459768
rect 316000 459756 316006 459808
rect 316586 459756 316592 459808
rect 316644 459796 316650 459808
rect 317322 459796 317328 459808
rect 316644 459768 317328 459796
rect 316644 459756 316650 459768
rect 317322 459756 317328 459768
rect 317380 459756 317386 459808
rect 318150 459756 318156 459808
rect 318208 459796 318214 459808
rect 318702 459796 318708 459808
rect 318208 459768 318708 459796
rect 318208 459756 318214 459768
rect 318702 459756 318708 459768
rect 318760 459756 318766 459808
rect 569218 459728 569224 459740
rect 287026 459700 569224 459728
rect 569218 459688 569224 459700
rect 569276 459688 569282 459740
rect 272334 459620 272340 459672
rect 272392 459660 272398 459672
rect 566458 459660 566464 459672
rect 272392 459632 566464 459660
rect 272392 459620 272398 459632
rect 566458 459620 566464 459632
rect 566516 459620 566522 459672
rect 267458 459552 267464 459604
rect 267516 459592 267522 459604
rect 562318 459592 562324 459604
rect 267516 459564 562324 459592
rect 267516 459552 267522 459564
rect 562318 459552 562324 459564
rect 562376 459552 562382 459604
rect 273990 458804 273996 458856
rect 274048 458844 274054 458856
rect 416038 458844 416044 458856
rect 274048 458816 416044 458844
rect 274048 458804 274054 458816
rect 416038 458804 416044 458816
rect 416096 458804 416102 458856
rect 231118 458736 231124 458788
rect 231176 458776 231182 458788
rect 374362 458776 374368 458788
rect 231176 458748 374368 458776
rect 231176 458736 231182 458748
rect 374362 458736 374368 458748
rect 374420 458736 374426 458788
rect 280062 458668 280068 458720
rect 280120 458708 280126 458720
rect 429838 458708 429844 458720
rect 280120 458680 429844 458708
rect 280120 458668 280126 458680
rect 429838 458668 429844 458680
rect 429896 458668 429902 458720
rect 222838 458600 222844 458652
rect 222896 458640 222902 458652
rect 375926 458640 375932 458652
rect 222896 458612 375932 458640
rect 222896 458600 222902 458612
rect 375926 458600 375932 458612
rect 375984 458600 375990 458652
rect 277026 458532 277032 458584
rect 277084 458572 277090 458584
rect 432598 458572 432604 458584
rect 277084 458544 432604 458572
rect 277084 458532 277090 458544
rect 432598 458532 432604 458544
rect 432656 458532 432662 458584
rect 232590 458464 232596 458516
rect 232648 458504 232654 458516
rect 391934 458504 391940 458516
rect 232648 458476 391940 458504
rect 232648 458464 232654 458476
rect 391934 458464 391940 458476
rect 391992 458464 391998 458516
rect 270402 458396 270408 458448
rect 270460 458436 270466 458448
rect 428550 458436 428556 458448
rect 270460 458408 428556 458436
rect 270460 458396 270466 458408
rect 428550 458396 428556 458408
rect 428608 458396 428614 458448
rect 228358 458328 228364 458380
rect 228416 458368 228422 458380
rect 407574 458368 407580 458380
rect 228416 458340 407580 458368
rect 228416 458328 228422 458340
rect 407574 458328 407580 458340
rect 407632 458328 407638 458380
rect 269022 458260 269028 458312
rect 269080 458300 269086 458312
rect 580258 458300 580264 458312
rect 269080 458272 580264 458300
rect 269080 458260 269086 458272
rect 580258 458260 580264 458272
rect 580316 458260 580322 458312
rect 3418 458192 3424 458244
rect 3476 458232 3482 458244
rect 373120 458232 373126 458244
rect 3476 458204 373126 458232
rect 3476 458192 3482 458204
rect 373120 458192 373126 458204
rect 373178 458192 373184 458244
rect 283466 457484 283472 457496
rect 283427 457456 283472 457484
rect 283466 457444 283472 457456
rect 283524 457444 283530 457496
rect 233878 457376 233884 457428
rect 233936 457416 233942 457428
rect 369854 457416 369860 457428
rect 233936 457388 369860 457416
rect 233936 457376 233942 457388
rect 369854 457376 369860 457388
rect 369912 457376 369918 457428
rect 377582 457416 377588 457428
rect 377543 457388 377588 457416
rect 377582 457376 377588 457388
rect 377640 457376 377646 457428
rect 379146 457416 379152 457428
rect 379107 457388 379152 457416
rect 379146 457376 379152 457388
rect 379204 457376 379210 457428
rect 380894 457416 380900 457428
rect 380855 457388 380900 457416
rect 380894 457376 380900 457388
rect 380952 457376 380958 457428
rect 278682 457308 278688 457360
rect 278740 457348 278746 457360
rect 418798 457348 418804 457360
rect 278740 457320 418804 457348
rect 278740 457308 278746 457320
rect 418798 457308 418804 457320
rect 418856 457308 418862 457360
rect 239214 457280 239220 457292
rect 239175 457252 239220 457280
rect 239214 457240 239220 457252
rect 239272 457240 239278 457292
rect 255038 457280 255044 457292
rect 254999 457252 255044 457280
rect 255038 457240 255044 457252
rect 255096 457240 255102 457292
rect 266078 457280 266084 457292
rect 266039 457252 266084 457280
rect 266078 457240 266084 457252
rect 266136 457240 266142 457292
rect 275554 457240 275560 457292
rect 275612 457280 275618 457292
rect 425698 457280 425704 457292
rect 275612 457252 425704 457280
rect 275612 457240 275618 457252
rect 425698 457240 425704 457252
rect 425756 457240 425762 457292
rect 226978 457172 226984 457224
rect 227036 457212 227042 457224
rect 379149 457215 379207 457221
rect 379149 457212 379161 457215
rect 227036 457184 379161 457212
rect 227036 457172 227042 457184
rect 379149 457181 379161 457184
rect 379195 457181 379207 457215
rect 379149 457175 379207 457181
rect 266081 457147 266139 457153
rect 266081 457113 266093 457147
rect 266127 457144 266139 457147
rect 421650 457144 421656 457156
rect 266127 457116 421656 457144
rect 266127 457113 266139 457116
rect 266081 457107 266139 457113
rect 421650 457104 421656 457116
rect 421708 457104 421714 457156
rect 224218 457036 224224 457088
rect 224276 457076 224282 457088
rect 380897 457079 380955 457085
rect 380897 457076 380909 457079
rect 224276 457048 380909 457076
rect 224276 457036 224282 457048
rect 380897 457045 380909 457048
rect 380943 457045 380955 457079
rect 380897 457039 380955 457045
rect 255041 457011 255099 457017
rect 255041 456977 255053 457011
rect 255087 457008 255099 457011
rect 417418 457008 417424 457020
rect 255087 456980 417424 457008
rect 255087 456977 255099 456980
rect 255041 456971 255099 456977
rect 417418 456968 417424 456980
rect 417476 456968 417482 457020
rect 239217 456943 239275 456949
rect 239217 456909 239229 456943
rect 239263 456940 239275 456943
rect 431218 456940 431224 456952
rect 239263 456912 431224 456940
rect 239263 456909 239275 456912
rect 239217 456903 239275 456909
rect 431218 456900 431224 456912
rect 431276 456900 431282 456952
rect 283469 456875 283527 456881
rect 283469 456841 283481 456875
rect 283515 456872 283527 456875
rect 579798 456872 579804 456884
rect 283515 456844 579804 456872
rect 283515 456841 283527 456844
rect 283469 456835 283527 456841
rect 579798 456832 579804 456844
rect 579856 456832 579862 456884
rect 4798 456764 4804 456816
rect 4856 456804 4862 456816
rect 377585 456807 377643 456813
rect 377585 456804 377597 456807
rect 4856 456776 377597 456804
rect 4856 456764 4862 456776
rect 377585 456773 377597 456776
rect 377631 456773 377643 456807
rect 377585 456767 377643 456773
rect 3326 449828 3332 449880
rect 3384 449868 3390 449880
rect 233878 449868 233884 449880
rect 3384 449840 233884 449868
rect 3384 449828 3390 449840
rect 233878 449828 233884 449840
rect 233936 449828 233942 449880
rect 429838 431876 429844 431928
rect 429896 431916 429902 431928
rect 580166 431916 580172 431928
rect 429896 431888 580172 431916
rect 429896 431876 429902 431888
rect 580166 431876 580172 431888
rect 580224 431876 580230 431928
rect 569218 419432 569224 419484
rect 569276 419472 569282 419484
rect 580166 419472 580172 419484
rect 569276 419444 580172 419472
rect 569276 419432 569282 419444
rect 580166 419432 580172 419444
rect 580224 419432 580230 419484
rect 3418 411204 3424 411256
rect 3476 411244 3482 411256
rect 222838 411244 222844 411256
rect 3476 411216 222844 411244
rect 3476 411204 3482 411216
rect 222838 411204 222844 411216
rect 222896 411204 222902 411256
rect 418798 405628 418804 405680
rect 418856 405668 418862 405680
rect 579614 405668 579620 405680
rect 418856 405640 579620 405668
rect 418856 405628 418862 405640
rect 579614 405628 579620 405640
rect 579672 405628 579678 405680
rect 3234 398760 3240 398812
rect 3292 398800 3298 398812
rect 231118 398800 231124 398812
rect 3292 398772 231124 398800
rect 3292 398760 3298 398772
rect 231118 398760 231124 398772
rect 231176 398760 231182 398812
rect 425698 379448 425704 379500
rect 425756 379488 425762 379500
rect 580166 379488 580172 379500
rect 425756 379460 580172 379488
rect 425756 379448 425762 379460
rect 580166 379448 580172 379460
rect 580224 379448 580230 379500
rect 2774 371424 2780 371476
rect 2832 371464 2838 371476
rect 4798 371464 4804 371476
rect 2832 371436 4804 371464
rect 2832 371424 2838 371436
rect 4798 371424 4804 371436
rect 4856 371424 4862 371476
rect 432598 365644 432604 365696
rect 432656 365684 432662 365696
rect 580166 365684 580172 365696
rect 432656 365656 580172 365684
rect 432656 365644 432662 365656
rect 580166 365644 580172 365656
rect 580224 365644 580230 365696
rect 3326 358708 3332 358760
rect 3384 358748 3390 358760
rect 224218 358748 224224 358760
rect 3384 358720 224224 358748
rect 3384 358708 3390 358720
rect 224218 358708 224224 358720
rect 224276 358708 224282 358760
rect 416038 353200 416044 353252
rect 416096 353240 416102 353252
rect 580166 353240 580172 353252
rect 416096 353212 580172 353240
rect 416096 353200 416102 353212
rect 580166 353200 580172 353212
rect 580224 353200 580230 353252
rect 3142 346332 3148 346384
rect 3200 346372 3206 346384
rect 226978 346372 226984 346384
rect 3200 346344 226984 346372
rect 3200 346332 3206 346344
rect 226978 346332 226984 346344
rect 227036 346332 227042 346384
rect 288452 336756 289952 336784
rect 220078 336676 220084 336728
rect 220136 336716 220142 336728
rect 288452 336716 288480 336756
rect 220136 336688 288480 336716
rect 220136 336676 220142 336688
rect 288526 336676 288532 336728
rect 288584 336716 288590 336728
rect 289814 336716 289820 336728
rect 288584 336688 289820 336716
rect 288584 336676 288590 336688
rect 289814 336676 289820 336688
rect 289872 336676 289878 336728
rect 289924 336716 289952 336756
rect 310514 336744 310520 336796
rect 310572 336784 310578 336796
rect 310790 336784 310796 336796
rect 310572 336756 310796 336784
rect 310572 336744 310578 336756
rect 310790 336744 310796 336756
rect 310848 336744 310854 336796
rect 289924 336688 290504 336716
rect 215938 336608 215944 336660
rect 215996 336648 216002 336660
rect 215996 336620 288388 336648
rect 215996 336608 216002 336620
rect 214558 336540 214564 336592
rect 214616 336580 214622 336592
rect 288253 336583 288311 336589
rect 288253 336580 288265 336583
rect 214616 336552 288265 336580
rect 214616 336540 214622 336552
rect 288253 336549 288265 336552
rect 288299 336549 288311 336583
rect 288360 336580 288388 336620
rect 288434 336608 288440 336660
rect 288492 336648 288498 336660
rect 289998 336648 290004 336660
rect 288492 336620 290004 336648
rect 288492 336608 288498 336620
rect 289998 336608 290004 336620
rect 290056 336608 290062 336660
rect 290476 336648 290504 336688
rect 291378 336676 291384 336728
rect 291436 336716 291442 336728
rect 292942 336716 292948 336728
rect 291436 336688 292948 336716
rect 291436 336676 291442 336688
rect 292942 336676 292948 336688
rect 293000 336676 293006 336728
rect 300486 336676 300492 336728
rect 300544 336716 300550 336728
rect 301314 336716 301320 336728
rect 300544 336688 301320 336716
rect 300544 336676 300550 336688
rect 301314 336676 301320 336688
rect 301372 336676 301378 336728
rect 304902 336676 304908 336728
rect 304960 336716 304966 336728
rect 328730 336716 328736 336728
rect 304960 336688 328736 336716
rect 304960 336676 304966 336688
rect 328730 336676 328736 336688
rect 328788 336676 328794 336728
rect 329190 336676 329196 336728
rect 329248 336716 329254 336728
rect 333974 336716 333980 336728
rect 329248 336688 333980 336716
rect 329248 336676 329254 336688
rect 333974 336676 333980 336688
rect 334032 336676 334038 336728
rect 339494 336676 339500 336728
rect 339552 336716 339558 336728
rect 339770 336716 339776 336728
rect 339552 336688 339776 336716
rect 339552 336676 339558 336688
rect 339770 336676 339776 336688
rect 339828 336676 339834 336728
rect 341610 336676 341616 336728
rect 341668 336716 341674 336728
rect 342070 336716 342076 336728
rect 341668 336688 342076 336716
rect 341668 336676 341674 336688
rect 342070 336676 342076 336688
rect 342128 336676 342134 336728
rect 343542 336676 343548 336728
rect 343600 336716 343606 336728
rect 344278 336716 344284 336728
rect 343600 336688 344284 336716
rect 343600 336676 343606 336688
rect 344278 336676 344284 336688
rect 344336 336676 344342 336728
rect 347038 336676 347044 336728
rect 347096 336716 347102 336728
rect 347682 336716 347688 336728
rect 347096 336688 347688 336716
rect 347096 336676 347102 336688
rect 347682 336676 347688 336688
rect 347740 336676 347746 336728
rect 348142 336676 348148 336728
rect 348200 336716 348206 336728
rect 349062 336716 349068 336728
rect 348200 336688 349068 336716
rect 348200 336676 348206 336688
rect 349062 336676 349068 336688
rect 349120 336676 349126 336728
rect 351086 336676 351092 336728
rect 351144 336716 351150 336728
rect 351822 336716 351828 336728
rect 351144 336688 351828 336716
rect 351144 336676 351150 336688
rect 351822 336676 351828 336688
rect 351880 336676 351886 336728
rect 352834 336676 352840 336728
rect 352892 336716 352898 336728
rect 353110 336716 353116 336728
rect 352892 336688 353116 336716
rect 352892 336676 352898 336688
rect 353110 336676 353116 336688
rect 353168 336676 353174 336728
rect 355686 336676 355692 336728
rect 355744 336716 355750 336728
rect 355962 336716 355968 336728
rect 355744 336688 355968 336716
rect 355744 336676 355750 336688
rect 355962 336676 355968 336688
rect 356020 336676 356026 336728
rect 357158 336676 357164 336728
rect 357216 336716 357222 336728
rect 357342 336716 357348 336728
rect 357216 336688 357348 336716
rect 357216 336676 357222 336688
rect 357342 336676 357348 336688
rect 357400 336676 357406 336728
rect 358354 336676 358360 336728
rect 358412 336716 358418 336728
rect 358630 336716 358636 336728
rect 358412 336688 358636 336716
rect 358412 336676 358418 336688
rect 358630 336676 358636 336688
rect 358688 336676 358694 336728
rect 360562 336676 360568 336728
rect 360620 336716 360626 336728
rect 361114 336716 361120 336728
rect 360620 336688 361120 336716
rect 360620 336676 360626 336688
rect 361114 336676 361120 336688
rect 361172 336676 361178 336728
rect 362586 336676 362592 336728
rect 362644 336716 362650 336728
rect 362862 336716 362868 336728
rect 362644 336688 362868 336716
rect 362644 336676 362650 336688
rect 362862 336676 362868 336688
rect 362920 336676 362926 336728
rect 363506 336676 363512 336728
rect 363564 336716 363570 336728
rect 364242 336716 364248 336728
rect 363564 336688 364248 336716
rect 363564 336676 363570 336688
rect 364242 336676 364248 336688
rect 364300 336676 364306 336728
rect 367462 336676 367468 336728
rect 367520 336716 367526 336728
rect 368290 336716 368296 336728
rect 367520 336688 368296 336716
rect 367520 336676 367526 336688
rect 368290 336676 368296 336688
rect 368348 336676 368354 336728
rect 368934 336676 368940 336728
rect 368992 336716 368998 336728
rect 369762 336716 369768 336728
rect 368992 336688 369768 336716
rect 368992 336676 368998 336688
rect 369762 336676 369768 336688
rect 369820 336676 369826 336728
rect 369854 336676 369860 336728
rect 369912 336716 369918 336728
rect 436094 336716 436100 336728
rect 369912 336688 436100 336716
rect 369912 336676 369918 336688
rect 436094 336676 436100 336688
rect 436152 336676 436158 336728
rect 294414 336648 294420 336660
rect 290476 336620 294420 336648
rect 294414 336608 294420 336620
rect 294472 336608 294478 336660
rect 296530 336608 296536 336660
rect 296588 336648 296594 336660
rect 296898 336648 296904 336660
rect 296588 336620 296904 336648
rect 296588 336608 296594 336620
rect 296898 336608 296904 336620
rect 296956 336608 296962 336660
rect 300762 336608 300768 336660
rect 300820 336648 300826 336660
rect 327534 336648 327540 336660
rect 300820 336620 327540 336648
rect 300820 336608 300826 336620
rect 327534 336608 327540 336620
rect 327592 336608 327598 336660
rect 355042 336608 355048 336660
rect 355100 336648 355106 336660
rect 355870 336648 355876 336660
rect 355100 336620 355876 336648
rect 355100 336608 355106 336620
rect 355870 336608 355876 336620
rect 355928 336608 355934 336660
rect 356808 336620 357848 336648
rect 292206 336580 292212 336592
rect 288360 336552 292212 336580
rect 288253 336543 288311 336549
rect 292206 336540 292212 336552
rect 292264 336540 292270 336592
rect 296622 336540 296628 336592
rect 296680 336580 296686 336592
rect 326154 336580 326160 336592
rect 296680 336552 326160 336580
rect 296680 336540 296686 336552
rect 326154 336540 326160 336552
rect 326212 336540 326218 336592
rect 327718 336540 327724 336592
rect 327776 336580 327782 336592
rect 328454 336580 328460 336592
rect 327776 336552 328460 336580
rect 327776 336540 327782 336552
rect 328454 336540 328460 336552
rect 328512 336540 328518 336592
rect 348418 336540 348424 336592
rect 348476 336580 348482 336592
rect 356808 336580 356836 336620
rect 348476 336552 356836 336580
rect 348476 336540 348482 336552
rect 356882 336540 356888 336592
rect 356940 336580 356946 336592
rect 357342 336580 357348 336592
rect 356940 336552 357348 336580
rect 356940 336540 356946 336552
rect 357342 336540 357348 336552
rect 357400 336540 357406 336592
rect 357820 336580 357848 336620
rect 357986 336608 357992 336660
rect 358044 336648 358050 336660
rect 358722 336648 358728 336660
rect 358044 336620 358728 336648
rect 358044 336608 358050 336620
rect 358722 336608 358728 336620
rect 358780 336608 358786 336660
rect 362034 336608 362040 336660
rect 362092 336648 362098 336660
rect 362678 336648 362684 336660
rect 362092 336620 362684 336648
rect 362092 336608 362098 336620
rect 362678 336608 362684 336620
rect 362736 336608 362742 336660
rect 366450 336608 366456 336660
rect 366508 336648 366514 336660
rect 367002 336648 367008 336660
rect 366508 336620 367008 336648
rect 366508 336608 366514 336620
rect 367002 336608 367008 336620
rect 367060 336608 367066 336660
rect 372246 336608 372252 336660
rect 372304 336648 372310 336660
rect 442994 336648 443000 336660
rect 372304 336620 443000 336648
rect 372304 336608 372310 336620
rect 442994 336608 443000 336620
rect 443052 336608 443058 336660
rect 363598 336580 363604 336592
rect 357820 336552 363604 336580
rect 363598 336540 363604 336552
rect 363656 336540 363662 336592
rect 373350 336540 373356 336592
rect 373408 336580 373414 336592
rect 373902 336580 373908 336592
rect 373408 336552 373908 336580
rect 373408 336540 373414 336552
rect 373902 336540 373908 336552
rect 373960 336540 373966 336592
rect 375926 336540 375932 336592
rect 375984 336580 375990 336592
rect 376662 336580 376668 336592
rect 375984 336552 376668 336580
rect 375984 336540 375990 336552
rect 376662 336540 376668 336552
rect 376720 336540 376726 336592
rect 377030 336540 377036 336592
rect 377088 336580 377094 336592
rect 377858 336580 377864 336592
rect 377088 336552 377864 336580
rect 377088 336540 377094 336552
rect 377858 336540 377864 336552
rect 377916 336540 377922 336592
rect 380250 336540 380256 336592
rect 380308 336580 380314 336592
rect 380710 336580 380716 336592
rect 380308 336552 380716 336580
rect 380308 336540 380314 336552
rect 380710 336540 380716 336552
rect 380768 336540 380774 336592
rect 381998 336540 382004 336592
rect 382056 336580 382062 336592
rect 382182 336580 382188 336592
rect 382056 336552 382188 336580
rect 382056 336540 382062 336552
rect 382182 336540 382188 336552
rect 382240 336540 382246 336592
rect 382277 336583 382335 336589
rect 382277 336549 382289 336583
rect 382323 336580 382335 336583
rect 449894 336580 449900 336592
rect 382323 336552 449900 336580
rect 382323 336549 382335 336552
rect 382277 336543 382335 336549
rect 449894 336540 449900 336552
rect 449952 336540 449958 336592
rect 209038 336472 209044 336524
rect 209096 336512 209102 336524
rect 296714 336512 296720 336524
rect 209096 336484 296720 336512
rect 209096 336472 209102 336484
rect 296714 336472 296720 336484
rect 296772 336472 296778 336524
rect 299382 336472 299388 336524
rect 299440 336512 299446 336524
rect 327074 336512 327080 336524
rect 299440 336484 327080 336512
rect 299440 336472 299446 336484
rect 327074 336472 327080 336484
rect 327132 336472 327138 336524
rect 347406 336472 347412 336524
rect 347464 336512 347470 336524
rect 358078 336512 358084 336524
rect 347464 336484 358084 336512
rect 347464 336472 347470 336484
rect 358078 336472 358084 336484
rect 358136 336472 358142 336524
rect 367830 336472 367836 336524
rect 367888 336512 367894 336524
rect 378781 336515 378839 336521
rect 378781 336512 378793 336515
rect 367888 336484 378793 336512
rect 367888 336472 367894 336484
rect 378781 336481 378793 336484
rect 378827 336481 378839 336515
rect 378781 336475 378839 336481
rect 379882 336472 379888 336524
rect 379940 336512 379946 336524
rect 380802 336512 380808 336524
rect 379940 336484 380808 336512
rect 379940 336472 379946 336484
rect 380802 336472 380808 336484
rect 380860 336472 380866 336524
rect 381354 336472 381360 336524
rect 381412 336512 381418 336524
rect 381906 336512 381912 336524
rect 381412 336484 381912 336512
rect 381412 336472 381418 336484
rect 381906 336472 381912 336484
rect 381964 336472 381970 336524
rect 456794 336512 456800 336524
rect 383626 336484 456800 336512
rect 125502 336404 125508 336456
rect 125560 336444 125566 336456
rect 273254 336444 273260 336456
rect 125560 336416 273260 336444
rect 125560 336404 125566 336416
rect 273254 336404 273260 336416
rect 273312 336404 273318 336456
rect 276014 336404 276020 336456
rect 276072 336444 276078 336456
rect 279050 336444 279056 336456
rect 276072 336416 279056 336444
rect 276072 336404 276078 336416
rect 279050 336404 279056 336416
rect 279108 336404 279114 336456
rect 282638 336404 282644 336456
rect 282696 336444 282702 336456
rect 283374 336444 283380 336456
rect 282696 336416 283380 336444
rect 282696 336404 282702 336416
rect 283374 336404 283380 336416
rect 283432 336404 283438 336456
rect 288253 336447 288311 336453
rect 288253 336413 288265 336447
rect 288299 336444 288311 336447
rect 293310 336444 293316 336456
rect 288299 336416 293316 336444
rect 288299 336413 288311 336416
rect 288253 336407 288311 336413
rect 293310 336404 293316 336416
rect 293368 336404 293374 336456
rect 293405 336447 293463 336453
rect 293405 336413 293417 336447
rect 293451 336444 293463 336447
rect 323578 336444 323584 336456
rect 293451 336416 323584 336444
rect 293451 336413 293463 336416
rect 293405 336407 293463 336413
rect 323578 336404 323584 336416
rect 323636 336404 323642 336456
rect 352190 336404 352196 336456
rect 352248 336444 352254 336456
rect 354585 336447 354643 336453
rect 354585 336444 354597 336447
rect 352248 336416 354597 336444
rect 352248 336404 352254 336416
rect 354585 336413 354597 336416
rect 354631 336413 354643 336447
rect 354585 336407 354643 336413
rect 369302 336404 369308 336456
rect 369360 336444 369366 336456
rect 378689 336447 378747 336453
rect 378689 336444 378701 336447
rect 369360 336416 378701 336444
rect 369360 336404 369366 336416
rect 378689 336413 378701 336416
rect 378735 336413 378747 336447
rect 383626 336444 383654 336484
rect 456794 336472 456800 336484
rect 456852 336472 456858 336524
rect 378689 336407 378747 336413
rect 381648 336416 383654 336444
rect 114462 336336 114468 336388
rect 114520 336376 114526 336388
rect 269942 336376 269948 336388
rect 114520 336348 269948 336376
rect 114520 336336 114526 336348
rect 269942 336336 269948 336348
rect 270000 336336 270006 336388
rect 277302 336336 277308 336388
rect 277360 336376 277366 336388
rect 319898 336376 319904 336388
rect 277360 336348 319904 336376
rect 277360 336336 277366 336348
rect 319898 336336 319904 336348
rect 319956 336336 319962 336388
rect 346670 336336 346676 336388
rect 346728 336376 346734 336388
rect 347590 336376 347596 336388
rect 346728 336348 347596 336376
rect 346728 336336 346734 336348
rect 347590 336336 347596 336348
rect 347648 336336 347654 336388
rect 354398 336336 354404 336388
rect 354456 336376 354462 336388
rect 370498 336376 370504 336388
rect 354456 336348 370504 336376
rect 354456 336336 354462 336348
rect 370498 336336 370504 336348
rect 370556 336336 370562 336388
rect 376570 336336 376576 336388
rect 376628 336376 376634 336388
rect 381648 336376 381676 336416
rect 383930 336404 383936 336456
rect 383988 336444 383994 336456
rect 384850 336444 384856 336456
rect 383988 336416 384856 336444
rect 383988 336404 383994 336416
rect 384850 336404 384856 336416
rect 384908 336404 384914 336456
rect 387242 336404 387248 336456
rect 387300 336444 387306 336456
rect 387702 336444 387708 336456
rect 387300 336416 387708 336444
rect 387300 336404 387306 336416
rect 387702 336404 387708 336416
rect 387760 336404 387766 336456
rect 388346 336404 388352 336456
rect 388404 336444 388410 336456
rect 389082 336444 389088 336456
rect 388404 336416 389088 336444
rect 388404 336404 388410 336416
rect 389082 336404 389088 336416
rect 389140 336404 389146 336456
rect 389450 336404 389456 336456
rect 389508 336444 389514 336456
rect 390186 336444 390192 336456
rect 389508 336416 390192 336444
rect 389508 336404 389514 336416
rect 390186 336404 390192 336416
rect 390244 336404 390250 336456
rect 392670 336404 392676 336456
rect 392728 336444 392734 336456
rect 393130 336444 393136 336456
rect 392728 336416 393136 336444
rect 392728 336404 392734 336416
rect 393130 336404 393136 336416
rect 393188 336404 393194 336456
rect 393225 336447 393283 336453
rect 393225 336413 393237 336447
rect 393271 336444 393283 336447
rect 465074 336444 465080 336456
rect 393271 336416 465080 336444
rect 393271 336413 393283 336416
rect 393225 336407 393283 336413
rect 465074 336404 465080 336416
rect 465132 336404 465138 336456
rect 376628 336348 381676 336376
rect 376628 336336 376634 336348
rect 381722 336336 381728 336388
rect 381780 336376 381786 336388
rect 468478 336376 468484 336388
rect 381780 336348 468484 336376
rect 381780 336336 381786 336348
rect 468478 336336 468484 336348
rect 468536 336336 468542 336388
rect 107562 336268 107568 336320
rect 107620 336308 107626 336320
rect 267826 336308 267832 336320
rect 107620 336280 267832 336308
rect 107620 336268 107626 336280
rect 267826 336268 267832 336280
rect 267884 336268 267890 336320
rect 277394 336268 277400 336320
rect 277452 336308 277458 336320
rect 279786 336308 279792 336320
rect 277452 336280 279792 336308
rect 277452 336268 277458 336280
rect 279786 336268 279792 336280
rect 279844 336268 279850 336320
rect 282178 336268 282184 336320
rect 282236 336308 282242 336320
rect 283098 336308 283104 336320
rect 282236 336280 283104 336308
rect 282236 336268 282242 336280
rect 283098 336268 283104 336280
rect 283156 336268 283162 336320
rect 283193 336311 283251 336317
rect 283193 336277 283205 336311
rect 283239 336308 283251 336311
rect 321554 336308 321560 336320
rect 283239 336280 321560 336308
rect 283239 336277 283251 336280
rect 283193 336271 283251 336277
rect 321554 336268 321560 336280
rect 321612 336268 321618 336320
rect 346302 336268 346308 336320
rect 346360 336308 346366 336320
rect 347130 336308 347136 336320
rect 346360 336280 347136 336308
rect 346360 336268 346366 336280
rect 347130 336268 347136 336280
rect 347188 336268 347194 336320
rect 348878 336268 348884 336320
rect 348936 336308 348942 336320
rect 367462 336308 367468 336320
rect 348936 336280 367468 336308
rect 348936 336268 348942 336280
rect 367462 336268 367468 336280
rect 367520 336268 367526 336320
rect 380986 336268 380992 336320
rect 381044 336308 381050 336320
rect 471974 336308 471980 336320
rect 381044 336280 471980 336308
rect 381044 336268 381050 336280
rect 471974 336268 471980 336280
rect 472032 336268 472038 336320
rect 57238 336200 57244 336252
rect 57296 336240 57302 336252
rect 251266 336240 251272 336252
rect 57296 336212 251272 336240
rect 57296 336200 57302 336212
rect 251266 336200 251272 336212
rect 251324 336200 251330 336252
rect 259454 336200 259460 336252
rect 259512 336240 259518 336252
rect 261478 336240 261484 336252
rect 259512 336212 261484 336240
rect 259512 336200 259518 336212
rect 261478 336200 261484 336212
rect 261536 336200 261542 336252
rect 264514 336200 264520 336252
rect 264572 336240 264578 336252
rect 265158 336240 265164 336252
rect 264572 336212 265164 336240
rect 264572 336200 264578 336212
rect 265158 336200 265164 336212
rect 265216 336200 265222 336252
rect 270034 336200 270040 336252
rect 270092 336240 270098 336252
rect 271874 336240 271880 336252
rect 270092 336212 271880 336240
rect 270092 336200 270098 336212
rect 271874 336200 271880 336212
rect 271932 336200 271938 336252
rect 274542 336200 274548 336252
rect 274600 336240 274606 336252
rect 319254 336240 319260 336252
rect 274600 336212 319260 336240
rect 274600 336200 274606 336212
rect 319254 336200 319260 336212
rect 319312 336200 319318 336252
rect 354030 336200 354036 336252
rect 354088 336240 354094 336252
rect 354490 336240 354496 336252
rect 354088 336212 354496 336240
rect 354088 336200 354094 336212
rect 354490 336200 354496 336212
rect 354548 336200 354554 336252
rect 354585 336243 354643 336249
rect 354585 336209 354597 336243
rect 354631 336240 354643 336243
rect 371786 336240 371792 336252
rect 354631 336212 371792 336240
rect 354631 336209 354643 336212
rect 354585 336203 354643 336209
rect 371786 336200 371792 336212
rect 371844 336200 371850 336252
rect 374454 336200 374460 336252
rect 374512 336240 374518 336252
rect 382277 336243 382335 336249
rect 382277 336240 382289 336243
rect 374512 336212 382289 336240
rect 374512 336200 374518 336212
rect 382277 336209 382289 336212
rect 382323 336209 382335 336243
rect 382277 336203 382335 336209
rect 383470 336200 383476 336252
rect 383528 336240 383534 336252
rect 475378 336240 475384 336252
rect 383528 336212 475384 336240
rect 383528 336200 383534 336212
rect 475378 336200 475384 336212
rect 475436 336200 475442 336252
rect 51718 336132 51724 336184
rect 51776 336172 51782 336184
rect 247954 336172 247960 336184
rect 51776 336144 247960 336172
rect 51776 336132 51782 336144
rect 247954 336132 247960 336144
rect 248012 336132 248018 336184
rect 267642 336132 267648 336184
rect 267700 336172 267706 336184
rect 317046 336172 317052 336184
rect 267700 336144 317052 336172
rect 267700 336132 267706 336144
rect 317046 336132 317052 336144
rect 317104 336132 317110 336184
rect 344094 336132 344100 336184
rect 344152 336172 344158 336184
rect 345658 336172 345664 336184
rect 344152 336144 345664 336172
rect 344152 336132 344158 336144
rect 345658 336132 345664 336144
rect 345716 336132 345722 336184
rect 351454 336132 351460 336184
rect 351512 336172 351518 336184
rect 375466 336172 375472 336184
rect 351512 336144 375472 336172
rect 351512 336132 351518 336144
rect 375466 336132 375472 336144
rect 375524 336132 375530 336184
rect 382458 336172 382464 336184
rect 378244 336144 382464 336172
rect 50338 336064 50344 336116
rect 50396 336104 50402 336116
rect 245838 336104 245844 336116
rect 50396 336076 245844 336104
rect 50396 336064 50402 336076
rect 245838 336064 245844 336076
rect 245896 336064 245902 336116
rect 270402 336064 270408 336116
rect 270460 336104 270466 336116
rect 318150 336104 318156 336116
rect 270460 336076 318156 336104
rect 270460 336064 270466 336076
rect 318150 336064 318156 336076
rect 318208 336064 318214 336116
rect 328362 336064 328368 336116
rect 328420 336104 328426 336116
rect 335998 336104 336004 336116
rect 328420 336076 336004 336104
rect 328420 336064 328426 336076
rect 335998 336064 336004 336076
rect 336056 336064 336062 336116
rect 353662 336064 353668 336116
rect 353720 336104 353726 336116
rect 378244 336104 378272 336144
rect 382458 336132 382464 336144
rect 382516 336132 382522 336184
rect 383194 336132 383200 336184
rect 383252 336172 383258 336184
rect 478874 336172 478880 336184
rect 383252 336144 478880 336172
rect 383252 336132 383258 336144
rect 478874 336132 478880 336144
rect 478932 336132 478938 336184
rect 353720 336076 378272 336104
rect 353720 336064 353726 336076
rect 378870 336064 378876 336116
rect 378928 336104 378934 336116
rect 393133 336107 393191 336113
rect 393133 336104 393145 336107
rect 378928 336076 393145 336104
rect 378928 336064 378934 336076
rect 393133 336073 393145 336076
rect 393179 336073 393191 336107
rect 393133 336067 393191 336073
rect 393222 336064 393228 336116
rect 393280 336104 393286 336116
rect 497458 336104 497464 336116
rect 393280 336076 497464 336104
rect 393280 336064 393286 336076
rect 497458 336064 497464 336076
rect 497516 336064 497522 336116
rect 35158 335996 35164 336048
rect 35216 336036 35222 336048
rect 243630 336036 243636 336048
rect 35216 336008 243636 336036
rect 35216 335996 35222 336008
rect 243630 335996 243636 336008
rect 243688 335996 243694 336048
rect 263502 335996 263508 336048
rect 263560 336036 263566 336048
rect 316034 336036 316040 336048
rect 263560 336008 316040 336036
rect 263560 335996 263566 336008
rect 316034 335996 316040 336008
rect 316092 335996 316098 336048
rect 316678 335996 316684 336048
rect 316736 336036 316742 336048
rect 327258 336036 327264 336048
rect 316736 336008 327264 336036
rect 316736 335996 316742 336008
rect 327258 335996 327264 336008
rect 327316 335996 327322 336048
rect 333238 335996 333244 336048
rect 333296 336036 333302 336048
rect 336734 336036 336740 336048
rect 333296 336008 336740 336036
rect 333296 335996 333302 336008
rect 336734 335996 336740 336008
rect 336792 335996 336798 336048
rect 344830 335996 344836 336048
rect 344888 336036 344894 336048
rect 348418 336036 348424 336048
rect 344888 336008 348424 336036
rect 344888 335996 344894 336008
rect 348418 335996 348424 336008
rect 348476 335996 348482 336048
rect 356514 335996 356520 336048
rect 356572 336036 356578 336048
rect 388438 336036 388444 336048
rect 356572 336008 388444 336036
rect 356572 335996 356578 336008
rect 388438 335996 388444 336008
rect 388496 335996 388502 336048
rect 391198 335996 391204 336048
rect 391256 336036 391262 336048
rect 504358 336036 504364 336048
rect 391256 336008 504364 336036
rect 391256 335996 391262 336008
rect 504358 335996 504364 336008
rect 504416 335996 504422 336048
rect 204898 335928 204904 335980
rect 204956 335968 204962 335980
rect 276842 335968 276848 335980
rect 204956 335940 276848 335968
rect 204956 335928 204962 335940
rect 276842 335928 276848 335940
rect 276900 335928 276906 335980
rect 281350 335928 281356 335980
rect 281408 335968 281414 335980
rect 283193 335971 283251 335977
rect 283193 335968 283205 335971
rect 281408 335940 283205 335968
rect 281408 335928 281414 335940
rect 283193 335937 283205 335940
rect 283239 335937 283251 335971
rect 283193 335931 283251 335937
rect 286410 335928 286416 335980
rect 286468 335968 286474 335980
rect 315206 335968 315212 335980
rect 286468 335940 315212 335968
rect 286468 335928 286474 335940
rect 315206 335928 315212 335940
rect 315264 335928 315270 335980
rect 335998 335928 336004 335980
rect 336056 335968 336062 335980
rect 337470 335968 337476 335980
rect 336056 335940 337476 335968
rect 336056 335928 336062 335940
rect 337470 335928 337476 335940
rect 337528 335928 337534 335980
rect 370406 335928 370412 335980
rect 370464 335968 370470 335980
rect 435358 335968 435364 335980
rect 370464 335940 435364 335968
rect 370464 335928 370470 335940
rect 435358 335928 435364 335940
rect 435416 335928 435422 335980
rect 224218 335860 224224 335912
rect 224276 335900 224282 335912
rect 291194 335900 291200 335912
rect 224276 335872 291200 335900
rect 224276 335860 224282 335872
rect 291194 335860 291200 335872
rect 291252 335860 291258 335912
rect 291930 335860 291936 335912
rect 291988 335900 291994 335912
rect 311894 335900 311900 335912
rect 291988 335872 311900 335900
rect 291988 335860 291994 335872
rect 311894 335860 311900 335872
rect 311952 335860 311958 335912
rect 366910 335860 366916 335912
rect 366968 335900 366974 335912
rect 366968 335872 372476 335900
rect 366968 335860 366974 335872
rect 233878 335792 233884 335844
rect 233936 335832 233942 335844
rect 300210 335832 300216 335844
rect 233936 335804 300216 335832
rect 233936 335792 233942 335804
rect 300210 335792 300216 335804
rect 300268 335792 300274 335844
rect 345566 335792 345572 335844
rect 345624 335832 345630 335844
rect 349798 335832 349804 335844
rect 345624 335804 349804 335832
rect 345624 335792 345630 335804
rect 349798 335792 349804 335804
rect 349856 335792 349862 335844
rect 359090 335792 359096 335844
rect 359148 335832 359154 335844
rect 360010 335832 360016 335844
rect 359148 335804 360016 335832
rect 359148 335792 359154 335804
rect 360010 335792 360016 335804
rect 360068 335792 360074 335844
rect 371878 335792 371884 335844
rect 371936 335832 371942 335844
rect 372338 335832 372344 335844
rect 371936 335804 372344 335832
rect 371936 335792 371942 335804
rect 372338 335792 372344 335804
rect 372396 335792 372402 335844
rect 372448 335832 372476 335872
rect 372982 335860 372988 335912
rect 373040 335900 373046 335912
rect 374638 335900 374644 335912
rect 373040 335872 374644 335900
rect 373040 335860 373046 335872
rect 374638 335860 374644 335872
rect 374696 335860 374702 335912
rect 378781 335903 378839 335909
rect 378781 335869 378793 335903
rect 378827 335900 378839 335903
rect 429194 335900 429200 335912
rect 378827 335872 429200 335900
rect 378827 335869 378839 335872
rect 378781 335863 378839 335869
rect 429194 335860 429200 335872
rect 429252 335860 429258 335912
rect 425698 335832 425704 335844
rect 372448 335804 425704 335832
rect 425698 335792 425704 335804
rect 425756 335792 425762 335844
rect 222838 335724 222844 335776
rect 222896 335764 222902 335776
rect 287790 335764 287796 335776
rect 222896 335736 287796 335764
rect 222896 335724 222902 335736
rect 287790 335724 287796 335736
rect 287848 335724 287854 335776
rect 289078 335724 289084 335776
rect 289136 335764 289142 335776
rect 312998 335764 313004 335776
rect 289136 335736 313004 335764
rect 289136 335724 289142 335736
rect 312998 335724 313004 335736
rect 313056 335724 313062 335776
rect 352558 335724 352564 335776
rect 352616 335764 352622 335776
rect 353202 335764 353208 335776
rect 352616 335736 353208 335764
rect 352616 335724 352622 335736
rect 353202 335724 353208 335736
rect 353260 335724 353266 335776
rect 378689 335767 378747 335773
rect 378689 335733 378701 335767
rect 378735 335764 378747 335767
rect 428458 335764 428464 335776
rect 378735 335736 428464 335764
rect 378735 335733 378747 335736
rect 378689 335727 378747 335733
rect 428458 335724 428464 335736
rect 428516 335724 428522 335776
rect 226978 335656 226984 335708
rect 227036 335696 227042 335708
rect 288894 335696 288900 335708
rect 227036 335668 288900 335696
rect 227036 335656 227042 335668
rect 288894 335656 288900 335668
rect 288952 335656 288958 335708
rect 295978 335656 295984 335708
rect 296036 335696 296042 335708
rect 314930 335696 314936 335708
rect 296036 335668 314936 335696
rect 296036 335656 296042 335668
rect 314930 335656 314936 335668
rect 314988 335656 314994 335708
rect 342714 335656 342720 335708
rect 342772 335696 342778 335708
rect 343358 335696 343364 335708
rect 342772 335668 343364 335696
rect 342772 335656 342778 335668
rect 343358 335656 343364 335668
rect 343416 335656 343422 335708
rect 349614 335656 349620 335708
rect 349672 335696 349678 335708
rect 353938 335696 353944 335708
rect 349672 335668 353944 335696
rect 349672 335656 349678 335668
rect 353938 335656 353944 335668
rect 353996 335656 354002 335708
rect 361206 335656 361212 335708
rect 361264 335696 361270 335708
rect 361482 335696 361488 335708
rect 361264 335668 361488 335696
rect 361264 335656 361270 335668
rect 361482 335656 361488 335668
rect 361540 335656 361546 335708
rect 366818 335656 366824 335708
rect 366876 335696 366882 335708
rect 425054 335696 425060 335708
rect 366876 335668 425060 335696
rect 366876 335656 366882 335668
rect 425054 335656 425060 335668
rect 425112 335656 425118 335708
rect 213178 335588 213184 335640
rect 213236 335628 213242 335640
rect 273898 335628 273904 335640
rect 213236 335600 273904 335628
rect 213236 335588 213242 335600
rect 273898 335588 273904 335600
rect 273956 335588 273962 335640
rect 288342 335588 288348 335640
rect 288400 335628 288406 335640
rect 293405 335631 293463 335637
rect 293405 335628 293417 335631
rect 288400 335600 293417 335628
rect 288400 335588 288406 335600
rect 293405 335597 293417 335600
rect 293451 335597 293463 335631
rect 293405 335591 293463 335597
rect 296438 335588 296444 335640
rect 296496 335628 296502 335640
rect 298094 335628 298100 335640
rect 296496 335600 298100 335628
rect 296496 335588 296502 335600
rect 298094 335588 298100 335600
rect 298152 335588 298158 335640
rect 366082 335588 366088 335640
rect 366140 335628 366146 335640
rect 413097 335631 413155 335637
rect 413097 335628 413109 335631
rect 366140 335600 413109 335628
rect 366140 335588 366146 335600
rect 413097 335597 413109 335600
rect 413143 335597 413155 335631
rect 413097 335591 413155 335597
rect 413186 335588 413192 335640
rect 413244 335628 413250 335640
rect 413830 335628 413836 335640
rect 413244 335600 413836 335628
rect 413244 335588 413250 335600
rect 413830 335588 413836 335600
rect 413888 335588 413894 335640
rect 414477 335631 414535 335637
rect 414477 335597 414489 335631
rect 414523 335628 414535 335631
rect 414753 335631 414811 335637
rect 414753 335628 414765 335631
rect 414523 335600 414765 335628
rect 414523 335597 414535 335600
rect 414477 335591 414535 335597
rect 414753 335597 414765 335600
rect 414799 335597 414811 335631
rect 414753 335591 414811 335597
rect 414842 335588 414848 335640
rect 414900 335628 414906 335640
rect 415118 335628 415124 335640
rect 414900 335600 415124 335628
rect 414900 335588 414906 335600
rect 415118 335588 415124 335600
rect 415176 335588 415182 335640
rect 415213 335631 415271 335637
rect 415213 335597 415225 335631
rect 415259 335628 415271 335631
rect 421558 335628 421564 335640
rect 415259 335600 421564 335628
rect 415259 335597 415271 335600
rect 415213 335591 415271 335597
rect 421558 335588 421564 335600
rect 421616 335588 421622 335640
rect 231118 335520 231124 335572
rect 231176 335560 231182 335572
rect 285674 335560 285680 335572
rect 231176 335532 285680 335560
rect 231176 335520 231182 335532
rect 285674 335520 285680 335532
rect 285732 335520 285738 335572
rect 341242 335520 341248 335572
rect 341300 335560 341306 335572
rect 342346 335560 342352 335572
rect 341300 335532 342352 335560
rect 341300 335520 341306 335532
rect 342346 335520 342352 335532
rect 342404 335520 342410 335572
rect 347498 335520 347504 335572
rect 347556 335560 347562 335572
rect 348510 335560 348516 335572
rect 347556 335532 348516 335560
rect 347556 335520 347562 335532
rect 348510 335520 348516 335532
rect 348568 335520 348574 335572
rect 364978 335520 364984 335572
rect 365036 335560 365042 335572
rect 414569 335563 414627 335569
rect 414569 335560 414581 335563
rect 365036 335532 414581 335560
rect 365036 335520 365042 335532
rect 414569 335529 414581 335532
rect 414615 335529 414627 335563
rect 414569 335523 414627 335529
rect 414658 335520 414664 335572
rect 414716 335560 414722 335572
rect 415302 335560 415308 335572
rect 414716 335532 415308 335560
rect 414716 335520 414722 335532
rect 415302 335520 415308 335532
rect 415360 335520 415366 335572
rect 232498 335452 232504 335504
rect 232556 335492 232562 335504
rect 282362 335492 282368 335504
rect 232556 335464 282368 335492
rect 232556 335452 232562 335464
rect 282362 335452 282368 335464
rect 282420 335452 282426 335504
rect 344462 335452 344468 335504
rect 344520 335492 344526 335504
rect 346946 335492 346952 335504
rect 344520 335464 346952 335492
rect 344520 335452 344526 335464
rect 346946 335452 346952 335464
rect 347004 335452 347010 335504
rect 363874 335452 363880 335504
rect 363932 335492 363938 335504
rect 416774 335492 416780 335504
rect 363932 335464 416780 335492
rect 363932 335452 363938 335464
rect 416774 335452 416780 335464
rect 416832 335452 416838 335504
rect 233970 335384 233976 335436
rect 234028 335424 234034 335436
rect 273530 335424 273536 335436
rect 234028 335396 273536 335424
rect 234028 335384 234034 335396
rect 273530 335384 273536 335396
rect 273588 335384 273594 335436
rect 341978 335384 341984 335436
rect 342036 335424 342042 335436
rect 345106 335424 345112 335436
rect 342036 335396 345112 335424
rect 342036 335384 342042 335396
rect 345106 335384 345112 335396
rect 345164 335384 345170 335436
rect 350074 335384 350080 335436
rect 350132 335424 350138 335436
rect 350350 335424 350356 335436
rect 350132 335396 350356 335424
rect 350132 335384 350138 335396
rect 350350 335384 350356 335396
rect 350408 335384 350414 335436
rect 364610 335384 364616 335436
rect 364668 335424 364674 335436
rect 418154 335424 418160 335436
rect 364668 335396 418160 335424
rect 364668 335384 364674 335396
rect 418154 335384 418160 335396
rect 418212 335384 418218 335436
rect 267734 335316 267740 335368
rect 267792 335356 267798 335368
rect 272794 335356 272800 335368
rect 267792 335328 272800 335356
rect 267792 335316 267798 335328
rect 272794 335316 272800 335328
rect 272852 335316 272858 335368
rect 274450 335316 274456 335368
rect 274508 335356 274514 335368
rect 278774 335356 278780 335368
rect 274508 335328 278780 335356
rect 274508 335316 274514 335328
rect 278774 335316 278780 335328
rect 278832 335316 278838 335368
rect 295426 335356 295432 335368
rect 292500 335328 295432 335356
rect 197262 335248 197268 335300
rect 197320 335288 197326 335300
rect 292500 335288 292528 335328
rect 295426 335316 295432 335328
rect 295484 335316 295490 335368
rect 332502 335316 332508 335368
rect 332560 335356 332566 335368
rect 337102 335356 337108 335368
rect 332560 335328 337108 335356
rect 332560 335316 332566 335328
rect 337102 335316 337108 335328
rect 337160 335316 337166 335368
rect 344922 335316 344928 335368
rect 344980 335356 344986 335368
rect 345750 335356 345756 335368
rect 344980 335328 345756 335356
rect 344980 335316 344986 335328
rect 345750 335316 345756 335328
rect 345808 335316 345814 335368
rect 355410 335316 355416 335368
rect 355468 335356 355474 335368
rect 382918 335356 382924 335368
rect 355468 335328 382924 335356
rect 355468 335316 355474 335328
rect 382918 335316 382924 335328
rect 382976 335316 382982 335368
rect 384666 335316 384672 335368
rect 384724 335356 384730 335368
rect 387153 335359 387211 335365
rect 387153 335356 387165 335359
rect 384724 335328 387165 335356
rect 384724 335316 384730 335328
rect 387153 335325 387165 335328
rect 387199 335325 387211 335359
rect 387153 335319 387211 335325
rect 388990 335316 388996 335368
rect 389048 335356 389054 335368
rect 393222 335356 393228 335368
rect 389048 335328 393228 335356
rect 389048 335316 389054 335328
rect 393222 335316 393228 335328
rect 393280 335316 393286 335368
rect 397822 335316 397828 335368
rect 397880 335356 397886 335368
rect 398558 335356 398564 335368
rect 397880 335328 398564 335356
rect 397880 335316 397886 335328
rect 398558 335316 398564 335328
rect 398616 335316 398622 335368
rect 402238 335316 402244 335368
rect 402296 335356 402302 335368
rect 402698 335356 402704 335368
rect 402296 335328 402704 335356
rect 402296 335316 402302 335328
rect 402698 335316 402704 335328
rect 402756 335316 402762 335368
rect 403986 335316 403992 335368
rect 404044 335356 404050 335368
rect 404262 335356 404268 335368
rect 404044 335328 404268 335356
rect 404044 335316 404050 335328
rect 404262 335316 404268 335328
rect 404320 335316 404326 335368
rect 405182 335316 405188 335368
rect 405240 335356 405246 335368
rect 405550 335356 405556 335368
rect 405240 335328 405556 335356
rect 405240 335316 405246 335328
rect 405550 335316 405556 335328
rect 405608 335316 405614 335368
rect 406562 335316 406568 335368
rect 406620 335356 406626 335368
rect 406838 335356 406844 335368
rect 406620 335328 406844 335356
rect 406620 335316 406626 335328
rect 406838 335316 406844 335328
rect 406896 335316 406902 335368
rect 407666 335316 407672 335368
rect 407724 335356 407730 335368
rect 408310 335356 408316 335368
rect 407724 335328 408316 335356
rect 407724 335316 407730 335328
rect 408310 335316 408316 335328
rect 408368 335316 408374 335368
rect 409506 335316 409512 335368
rect 409564 335356 409570 335368
rect 409782 335356 409788 335368
rect 409564 335328 409788 335356
rect 409564 335316 409570 335328
rect 409782 335316 409788 335328
rect 409840 335316 409846 335368
rect 410702 335316 410708 335368
rect 410760 335356 410766 335368
rect 411070 335356 411076 335368
rect 410760 335328 411076 335356
rect 410760 335316 410766 335328
rect 411070 335316 411076 335328
rect 411128 335316 411134 335368
rect 412082 335316 412088 335368
rect 412140 335356 412146 335368
rect 412358 335356 412364 335368
rect 412140 335328 412364 335356
rect 412140 335316 412146 335328
rect 412358 335316 412364 335328
rect 412416 335316 412422 335368
rect 413097 335359 413155 335365
rect 413097 335325 413109 335359
rect 413143 335356 413155 335359
rect 414477 335359 414535 335365
rect 414477 335356 414489 335359
rect 413143 335328 414489 335356
rect 413143 335325 413155 335328
rect 413097 335319 413155 335325
rect 414477 335325 414489 335328
rect 414523 335325 414535 335359
rect 414477 335319 414535 335325
rect 414569 335359 414627 335365
rect 414569 335325 414581 335359
rect 414615 335356 414627 335359
rect 418798 335356 418804 335368
rect 414615 335328 418804 335356
rect 414615 335325 414627 335328
rect 414569 335319 414627 335325
rect 418798 335316 418804 335328
rect 418856 335316 418862 335368
rect 197320 335260 292528 335288
rect 197320 335248 197326 335260
rect 373718 335248 373724 335300
rect 373776 335288 373782 335300
rect 448514 335288 448520 335300
rect 373776 335260 448520 335288
rect 373776 335248 373782 335260
rect 448514 335248 448520 335260
rect 448572 335248 448578 335300
rect 179322 335180 179328 335232
rect 179380 335220 179386 335232
rect 288434 335220 288440 335232
rect 179380 335192 288440 335220
rect 179380 335180 179386 335192
rect 288434 335180 288440 335192
rect 288492 335180 288498 335232
rect 387153 335223 387211 335229
rect 387153 335189 387165 335223
rect 387199 335220 387211 335223
rect 483014 335220 483020 335232
rect 387199 335192 483020 335220
rect 387199 335189 387211 335192
rect 387153 335183 387211 335189
rect 483014 335180 483020 335192
rect 483072 335180 483078 335232
rect 169662 335112 169668 335164
rect 169720 335152 169726 335164
rect 286686 335152 286692 335164
rect 169720 335124 286692 335152
rect 169720 335112 169726 335124
rect 286686 335112 286692 335124
rect 286744 335112 286750 335164
rect 384298 335112 384304 335164
rect 384356 335152 384362 335164
rect 481634 335152 481640 335164
rect 384356 335124 481640 335152
rect 384356 335112 384362 335124
rect 481634 335112 481640 335124
rect 481692 335112 481698 335164
rect 161382 335044 161388 335096
rect 161440 335084 161446 335096
rect 284478 335084 284484 335096
rect 161440 335056 284484 335084
rect 161440 335044 161446 335056
rect 284478 335044 284484 335056
rect 284536 335044 284542 335096
rect 391934 335044 391940 335096
rect 391992 335084 391998 335096
rect 490006 335084 490012 335096
rect 391992 335056 490012 335084
rect 391992 335044 391998 335056
rect 490006 335044 490012 335056
rect 490064 335044 490070 335096
rect 144822 334976 144828 335028
rect 144880 335016 144886 335028
rect 276014 335016 276020 335028
rect 144880 334988 276020 335016
rect 144880 334976 144886 334988
rect 276014 334976 276020 334988
rect 276072 334976 276078 335028
rect 390094 334976 390100 335028
rect 390152 335016 390158 335028
rect 500954 335016 500960 335028
rect 390152 334988 500960 335016
rect 390152 334976 390158 334988
rect 500954 334976 500960 334988
rect 501012 334976 501018 335028
rect 147582 334908 147588 334960
rect 147640 334948 147646 334960
rect 280246 334948 280252 334960
rect 147640 334920 280252 334948
rect 147640 334908 147646 334920
rect 280246 334908 280252 334920
rect 280304 334908 280310 334960
rect 392302 334908 392308 334960
rect 392360 334948 392366 334960
rect 507854 334948 507860 334960
rect 392360 334920 507860 334948
rect 392360 334908 392366 334920
rect 507854 334908 507860 334920
rect 507912 334908 507918 334960
rect 140682 334840 140688 334892
rect 140740 334880 140746 334892
rect 277946 334880 277952 334892
rect 140740 334852 277952 334880
rect 140740 334840 140746 334852
rect 277946 334840 277952 334852
rect 278004 334840 278010 334892
rect 393774 334840 393780 334892
rect 393832 334880 393838 334892
rect 512638 334880 512644 334892
rect 393832 334852 512644 334880
rect 393832 334840 393838 334852
rect 512638 334840 512644 334852
rect 512696 334840 512702 334892
rect 87598 334772 87604 334824
rect 87656 334812 87662 334824
rect 260926 334812 260932 334824
rect 87656 334784 260932 334812
rect 87656 334772 87662 334784
rect 260926 334772 260932 334784
rect 260984 334772 260990 334824
rect 398190 334772 398196 334824
rect 398248 334812 398254 334824
rect 526438 334812 526444 334824
rect 398248 334784 526444 334812
rect 398248 334772 398254 334784
rect 526438 334772 526444 334784
rect 526496 334772 526502 334824
rect 86862 334704 86868 334756
rect 86920 334744 86926 334756
rect 259454 334744 259460 334756
rect 86920 334716 259460 334744
rect 86920 334704 86926 334716
rect 259454 334704 259460 334716
rect 259512 334704 259518 334756
rect 397086 334704 397092 334756
rect 397144 334744 397150 334756
rect 522298 334744 522304 334756
rect 397144 334716 522304 334744
rect 397144 334704 397150 334716
rect 522298 334704 522304 334716
rect 522356 334704 522362 334756
rect 29638 334636 29644 334688
rect 29696 334676 29702 334688
rect 243262 334676 243268 334688
rect 29696 334648 243268 334676
rect 29696 334636 29702 334648
rect 243262 334636 243268 334648
rect 243320 334636 243326 334688
rect 398466 334636 398472 334688
rect 398524 334676 398530 334688
rect 528554 334676 528560 334688
rect 398524 334648 528560 334676
rect 398524 334636 398530 334648
rect 528554 334636 528560 334648
rect 528612 334636 528618 334688
rect 22738 334568 22744 334620
rect 22796 334608 22802 334620
rect 238846 334608 238852 334620
rect 22796 334580 238852 334608
rect 22796 334568 22802 334580
rect 238846 334568 238852 334580
rect 238904 334568 238910 334620
rect 402514 334568 402520 334620
rect 402572 334608 402578 334620
rect 540238 334608 540244 334620
rect 402572 334580 540244 334608
rect 402572 334568 402578 334580
rect 540238 334568 540244 334580
rect 540296 334568 540302 334620
rect 202782 334500 202788 334552
rect 202840 334540 202846 334552
rect 296530 334540 296536 334552
rect 202840 334512 296536 334540
rect 202840 334500 202846 334512
rect 296530 334500 296536 334512
rect 296588 334500 296594 334552
rect 371510 334500 371516 334552
rect 371568 334540 371574 334552
rect 440326 334540 440332 334552
rect 371568 334512 440332 334540
rect 371568 334500 371574 334512
rect 440326 334500 440332 334512
rect 440384 334500 440390 334552
rect 216582 334432 216588 334484
rect 216640 334472 216646 334484
rect 300486 334472 300492 334484
rect 216640 334444 300492 334472
rect 216640 334432 216646 334444
rect 300486 334432 300492 334444
rect 300544 334432 300550 334484
rect 368106 334432 368112 334484
rect 368164 334472 368170 334484
rect 430574 334472 430580 334484
rect 368164 334444 430580 334472
rect 368164 334432 368170 334444
rect 430574 334432 430580 334444
rect 430632 334432 430638 334484
rect 223482 334364 223488 334416
rect 223540 334404 223546 334416
rect 303614 334404 303620 334416
rect 223540 334376 303620 334404
rect 223540 334364 223546 334376
rect 303614 334364 303620 334376
rect 303672 334364 303678 334416
rect 205542 333888 205548 333940
rect 205600 333928 205606 333940
rect 296438 333928 296444 333940
rect 205600 333900 296444 333928
rect 205600 333888 205606 333900
rect 296438 333888 296444 333900
rect 296496 333888 296502 333940
rect 374638 333888 374644 333940
rect 374696 333928 374702 333940
rect 445754 333928 445760 333940
rect 374696 333900 445760 333928
rect 374696 333888 374702 333900
rect 445754 333888 445760 333900
rect 445812 333888 445818 333940
rect 198642 333820 198648 333872
rect 198700 333860 198706 333872
rect 295794 333860 295800 333872
rect 198700 333832 295800 333860
rect 198700 333820 198706 333832
rect 295794 333820 295800 333832
rect 295852 333820 295858 333872
rect 373810 333820 373816 333872
rect 373868 333860 373874 333872
rect 448606 333860 448612 333872
rect 373868 333832 448612 333860
rect 373868 333820 373874 333832
rect 448606 333820 448612 333832
rect 448664 333820 448670 333872
rect 177942 333752 177948 333804
rect 178000 333792 178006 333804
rect 288526 333792 288532 333804
rect 178000 333764 288532 333792
rect 178000 333752 178006 333764
rect 288526 333752 288532 333764
rect 288584 333752 288590 333804
rect 377398 333752 377404 333804
rect 377456 333792 377462 333804
rect 459554 333792 459560 333804
rect 377456 333764 459560 333792
rect 377456 333752 377462 333764
rect 459554 333752 459560 333764
rect 459612 333752 459618 333804
rect 162762 333684 162768 333736
rect 162820 333724 162826 333736
rect 284846 333724 284852 333736
rect 162820 333696 284852 333724
rect 162820 333684 162826 333696
rect 284846 333684 284852 333696
rect 284904 333684 284910 333736
rect 380894 333684 380900 333736
rect 380952 333724 380958 333736
rect 470594 333724 470600 333736
rect 380952 333696 470600 333724
rect 380952 333684 380958 333696
rect 470594 333684 470600 333696
rect 470652 333684 470658 333736
rect 158622 333616 158628 333668
rect 158680 333656 158686 333668
rect 282638 333656 282644 333668
rect 158680 333628 282644 333656
rect 158680 333616 158686 333628
rect 282638 333616 282644 333628
rect 282696 333616 282702 333668
rect 387610 333616 387616 333668
rect 387668 333656 387674 333668
rect 492674 333656 492680 333668
rect 387668 333628 492680 333656
rect 387668 333616 387674 333628
rect 492674 333616 492680 333628
rect 492732 333616 492738 333668
rect 151722 333548 151728 333600
rect 151780 333588 151786 333600
rect 281442 333588 281448 333600
rect 151780 333560 281448 333588
rect 151780 333548 151786 333560
rect 281442 333548 281448 333560
rect 281500 333548 281506 333600
rect 390922 333548 390928 333600
rect 390980 333588 390986 333600
rect 502978 333588 502984 333600
rect 390980 333560 502984 333588
rect 390980 333548 390986 333560
rect 502978 333548 502984 333560
rect 503036 333548 503042 333600
rect 93118 333480 93124 333532
rect 93176 333520 93182 333532
rect 262950 333520 262956 333532
rect 93176 333492 262956 333520
rect 93176 333480 93182 333492
rect 262950 333480 262956 333492
rect 263008 333480 263014 333532
rect 394602 333480 394608 333532
rect 394660 333520 394666 333532
rect 515398 333520 515404 333532
rect 394660 333492 515404 333520
rect 394660 333480 394666 333492
rect 515398 333480 515404 333492
rect 515456 333480 515462 333532
rect 88978 333412 88984 333464
rect 89036 333452 89042 333464
rect 261938 333452 261944 333464
rect 89036 333424 261944 333452
rect 89036 333412 89042 333424
rect 261938 333412 261944 333424
rect 261996 333412 262002 333464
rect 395890 333412 395896 333464
rect 395948 333452 395954 333464
rect 520274 333452 520280 333464
rect 395948 333424 520280 333452
rect 395948 333412 395954 333424
rect 520274 333412 520280 333424
rect 520332 333412 520338 333464
rect 84102 333344 84108 333396
rect 84160 333384 84166 333396
rect 260374 333384 260380 333396
rect 84160 333356 260380 333384
rect 84160 333344 84166 333356
rect 260374 333344 260380 333356
rect 260432 333344 260438 333396
rect 400122 333344 400128 333396
rect 400180 333384 400186 333396
rect 407853 333387 407911 333393
rect 400180 333356 407804 333384
rect 400180 333344 400186 333356
rect 54478 333276 54484 333328
rect 54536 333316 54542 333328
rect 247586 333316 247592 333328
rect 54536 333288 247592 333316
rect 54536 333276 54542 333288
rect 247586 333276 247592 333288
rect 247644 333276 247650 333328
rect 407776 333316 407804 333356
rect 407853 333353 407865 333387
rect 407899 333384 407911 333387
rect 530578 333384 530584 333396
rect 407899 333356 530584 333384
rect 407899 333353 407911 333356
rect 407853 333347 407911 333353
rect 530578 333344 530584 333356
rect 530636 333344 530642 333396
rect 533338 333316 533344 333328
rect 407776 333288 533344 333316
rect 533338 333276 533344 333288
rect 533396 333276 533402 333328
rect 39298 333208 39304 333260
rect 39356 333248 39362 333260
rect 241882 333248 241888 333260
rect 39356 333220 241888 333248
rect 39356 333208 39362 333220
rect 241882 333208 241888 333220
rect 241940 333208 241946 333260
rect 401502 333208 401508 333260
rect 401560 333248 401566 333260
rect 538214 333248 538220 333260
rect 401560 333220 538220 333248
rect 401560 333208 401566 333220
rect 538214 333208 538220 333220
rect 538272 333208 538278 333260
rect 209682 333140 209688 333192
rect 209740 333180 209746 333192
rect 299106 333180 299112 333192
rect 209740 333152 299112 333180
rect 209740 333140 209746 333152
rect 299106 333140 299112 333152
rect 299164 333140 299170 333192
rect 399294 333140 399300 333192
rect 399352 333180 399358 333192
rect 407853 333183 407911 333189
rect 407853 333180 407865 333183
rect 399352 333152 407865 333180
rect 399352 333140 399358 333152
rect 407853 333149 407865 333152
rect 407899 333149 407911 333183
rect 407853 333143 407911 333149
rect 227622 333072 227628 333124
rect 227680 333112 227686 333124
rect 304626 333112 304632 333124
rect 227680 333084 304632 333112
rect 227680 333072 227686 333084
rect 304626 333072 304632 333084
rect 304684 333072 304690 333124
rect 219250 332528 219256 332580
rect 219308 332568 219314 332580
rect 302418 332568 302424 332580
rect 219308 332540 302424 332568
rect 219308 332528 219314 332540
rect 302418 332528 302424 332540
rect 302476 332528 302482 332580
rect 188982 332460 188988 332512
rect 189040 332500 189046 332512
rect 291378 332500 291384 332512
rect 189040 332472 291384 332500
rect 189040 332460 189046 332472
rect 291378 332460 291384 332472
rect 291436 332460 291442 332512
rect 182082 332392 182088 332444
rect 182140 332432 182146 332444
rect 290826 332432 290832 332444
rect 182140 332404 290832 332432
rect 182140 332392 182146 332404
rect 290826 332392 290832 332404
rect 290884 332392 290890 332444
rect 375190 332392 375196 332444
rect 375248 332432 375254 332444
rect 452654 332432 452660 332444
rect 375248 332404 452660 332432
rect 375248 332392 375254 332404
rect 452654 332392 452660 332404
rect 452712 332392 452718 332444
rect 175182 332324 175188 332376
rect 175240 332364 175246 332376
rect 288618 332364 288624 332376
rect 175240 332336 288624 332364
rect 175240 332324 175246 332336
rect 288618 332324 288624 332336
rect 288676 332324 288682 332376
rect 376202 332324 376208 332376
rect 376260 332364 376266 332376
rect 456886 332364 456892 332376
rect 376260 332336 456892 332364
rect 376260 332324 376266 332336
rect 456886 332324 456892 332336
rect 456944 332324 456950 332376
rect 171042 332256 171048 332308
rect 171100 332296 171106 332308
rect 287422 332296 287428 332308
rect 171100 332268 287428 332296
rect 171100 332256 171106 332268
rect 287422 332256 287428 332268
rect 287480 332256 287486 332308
rect 378502 332256 378508 332308
rect 378560 332296 378566 332308
rect 463694 332296 463700 332308
rect 378560 332268 463700 332296
rect 378560 332256 378566 332268
rect 463694 332256 463700 332268
rect 463752 332256 463758 332308
rect 143442 332188 143448 332240
rect 143500 332228 143506 332240
rect 274450 332228 274456 332240
rect 143500 332200 274456 332228
rect 143500 332188 143506 332200
rect 274450 332188 274456 332200
rect 274508 332188 274514 332240
rect 379422 332188 379428 332240
rect 379480 332228 379486 332240
rect 466454 332228 466460 332240
rect 379480 332200 466460 332228
rect 379480 332188 379486 332200
rect 466454 332188 466460 332200
rect 466512 332188 466518 332240
rect 104158 332120 104164 332172
rect 104216 332160 104222 332172
rect 266354 332160 266360 332172
rect 104216 332132 266360 332160
rect 104216 332120 104222 332132
rect 266354 332120 266360 332132
rect 266412 332120 266418 332172
rect 382826 332120 382832 332172
rect 382884 332160 382890 332172
rect 477494 332160 477500 332172
rect 382884 332132 477500 332160
rect 382884 332120 382890 332132
rect 477494 332120 477500 332132
rect 477552 332120 477558 332172
rect 99282 332052 99288 332104
rect 99340 332092 99346 332104
rect 264514 332092 264520 332104
rect 99340 332064 264520 332092
rect 99340 332052 99346 332064
rect 264514 332052 264520 332064
rect 264572 332052 264578 332104
rect 385310 332052 385316 332104
rect 385368 332092 385374 332104
rect 485774 332092 485780 332104
rect 385368 332064 485780 332092
rect 385368 332052 385374 332064
rect 485774 332052 485780 332064
rect 485832 332052 485838 332104
rect 95142 331984 95148 332036
rect 95200 332024 95206 332036
rect 264054 332024 264060 332036
rect 95200 331996 264060 332024
rect 95200 331984 95206 331996
rect 264054 331984 264060 331996
rect 264112 331984 264118 332036
rect 388714 331984 388720 332036
rect 388772 332024 388778 332036
rect 496814 332024 496820 332036
rect 388772 331996 496820 332024
rect 388772 331984 388778 331996
rect 496814 331984 496820 331996
rect 496872 331984 496878 332036
rect 68278 331916 68284 331968
rect 68336 331956 68342 331968
rect 250162 331956 250168 331968
rect 68336 331928 250168 331956
rect 68336 331916 68342 331928
rect 250162 331916 250168 331928
rect 250220 331916 250226 331968
rect 391842 331916 391848 331968
rect 391900 331956 391906 331968
rect 506474 331956 506480 331968
rect 391900 331928 506480 331956
rect 391900 331916 391906 331928
rect 506474 331916 506480 331928
rect 506532 331916 506538 331968
rect 33778 331848 33784 331900
rect 33836 331888 33842 331900
rect 244458 331888 244464 331900
rect 33836 331860 244464 331888
rect 33836 331848 33842 331860
rect 244458 331848 244464 331860
rect 244516 331848 244522 331900
rect 396350 331848 396356 331900
rect 396408 331888 396414 331900
rect 519538 331888 519544 331900
rect 396408 331860 519544 331888
rect 396408 331848 396414 331860
rect 519538 331848 519544 331860
rect 519596 331848 519602 331900
rect 153102 330964 153108 331016
rect 153160 331004 153166 331016
rect 281994 331004 282000 331016
rect 153160 330976 282000 331004
rect 153160 330964 153166 330976
rect 281994 330964 282000 330976
rect 282052 330964 282058 331016
rect 146202 330896 146208 330948
rect 146260 330936 146266 330948
rect 277394 330936 277400 330948
rect 146260 330908 277400 330936
rect 146260 330896 146266 330908
rect 277394 330896 277400 330908
rect 277452 330896 277458 330948
rect 117222 330828 117228 330880
rect 117280 330868 117286 330880
rect 270862 330868 270868 330880
rect 117280 330840 270868 330868
rect 117280 330828 117286 330840
rect 270862 330828 270868 330840
rect 270920 330828 270926 330880
rect 399662 330828 399668 330880
rect 399720 330868 399726 330880
rect 485038 330868 485044 330880
rect 399720 330840 485044 330868
rect 399720 330828 399726 330840
rect 485038 330828 485044 330840
rect 485096 330828 485102 330880
rect 111058 330760 111064 330812
rect 111116 330800 111122 330812
rect 268470 330800 268476 330812
rect 111116 330772 268476 330800
rect 111116 330760 111122 330772
rect 268470 330760 268476 330772
rect 268528 330760 268534 330812
rect 324406 330760 324412 330812
rect 324464 330760 324470 330812
rect 386322 330760 386328 330812
rect 386380 330800 386386 330812
rect 489178 330800 489184 330812
rect 386380 330772 489184 330800
rect 386380 330760 386386 330772
rect 489178 330760 489184 330772
rect 489236 330760 489242 330812
rect 106182 330692 106188 330744
rect 106240 330732 106246 330744
rect 267366 330732 267372 330744
rect 106240 330704 267372 330732
rect 106240 330692 106246 330704
rect 267366 330692 267372 330704
rect 267424 330692 267430 330744
rect 81342 330624 81348 330676
rect 81400 330664 81406 330676
rect 259638 330664 259644 330676
rect 81400 330636 259644 330664
rect 81400 330624 81406 330636
rect 259638 330624 259644 330636
rect 259696 330624 259702 330676
rect 324424 330608 324452 330760
rect 389818 330692 389824 330744
rect 389876 330732 389882 330744
rect 499574 330732 499580 330744
rect 389876 330704 499580 330732
rect 389876 330692 389882 330704
rect 499574 330692 499580 330704
rect 499632 330692 499638 330744
rect 392854 330624 392860 330676
rect 392912 330664 392918 330676
rect 510614 330664 510620 330676
rect 392912 330636 510620 330664
rect 392912 330624 392918 330636
rect 510614 330624 510620 330636
rect 510672 330624 510678 330676
rect 58618 330556 58624 330608
rect 58676 330596 58682 330608
rect 248690 330596 248696 330608
rect 58676 330568 248696 330596
rect 58676 330556 58682 330568
rect 248690 330556 248696 330568
rect 248748 330556 248754 330608
rect 324406 330556 324412 330608
rect 324464 330556 324470 330608
rect 394142 330556 394148 330608
rect 394200 330596 394206 330608
rect 514754 330596 514760 330608
rect 394200 330568 514760 330596
rect 394200 330556 394206 330568
rect 514754 330556 514760 330568
rect 514812 330556 514818 330608
rect 36538 330488 36544 330540
rect 36596 330528 36602 330540
rect 36596 330500 238754 330528
rect 36596 330488 36602 330500
rect 234798 330420 234804 330472
rect 234856 330460 234862 330472
rect 235534 330460 235540 330472
rect 234856 330432 235540 330460
rect 234856 330420 234862 330432
rect 235534 330420 235540 330432
rect 235592 330420 235598 330472
rect 236086 330420 236092 330472
rect 236144 330460 236150 330472
rect 237006 330460 237012 330472
rect 236144 330432 237012 330460
rect 236144 330420 236150 330432
rect 237006 330420 237012 330432
rect 237064 330420 237070 330472
rect 237374 330420 237380 330472
rect 237432 330460 237438 330472
rect 238478 330460 238484 330472
rect 237432 330432 238484 330460
rect 237432 330420 237438 330432
rect 238478 330420 238484 330432
rect 238536 330420 238542 330472
rect 238726 330460 238754 330500
rect 241606 330488 241612 330540
rect 241664 330528 241670 330540
rect 242526 330528 242532 330540
rect 241664 330500 242532 330528
rect 241664 330488 241670 330500
rect 242526 330488 242532 330500
rect 242584 330488 242590 330540
rect 244366 330488 244372 330540
rect 244424 330528 244430 330540
rect 245102 330528 245108 330540
rect 244424 330500 245108 330528
rect 244424 330488 244430 330500
rect 245102 330488 245108 330500
rect 245160 330488 245166 330540
rect 247126 330488 247132 330540
rect 247184 330528 247190 330540
rect 247310 330528 247316 330540
rect 247184 330500 247316 330528
rect 247184 330488 247190 330500
rect 247310 330488 247316 330500
rect 247368 330488 247374 330540
rect 248506 330488 248512 330540
rect 248564 330528 248570 330540
rect 249426 330528 249432 330540
rect 248564 330500 249432 330528
rect 248564 330488 248570 330500
rect 249426 330488 249432 330500
rect 249484 330488 249490 330540
rect 249886 330488 249892 330540
rect 249944 330528 249950 330540
rect 250898 330528 250904 330540
rect 249944 330500 250904 330528
rect 249944 330488 249950 330500
rect 250898 330488 250904 330500
rect 250956 330488 250962 330540
rect 251266 330488 251272 330540
rect 251324 330528 251330 330540
rect 252002 330528 252008 330540
rect 251324 330500 252008 330528
rect 251324 330488 251330 330500
rect 252002 330488 252008 330500
rect 252060 330488 252066 330540
rect 253934 330488 253940 330540
rect 253992 330528 253998 330540
rect 254578 330528 254584 330540
rect 253992 330500 254584 330528
rect 253992 330488 253998 330500
rect 254578 330488 254584 330500
rect 254636 330488 254642 330540
rect 255406 330488 255412 330540
rect 255464 330528 255470 330540
rect 256050 330528 256056 330540
rect 255464 330500 256056 330528
rect 255464 330488 255470 330500
rect 256050 330488 256056 330500
rect 256108 330488 256114 330540
rect 258166 330488 258172 330540
rect 258224 330528 258230 330540
rect 258994 330528 259000 330540
rect 258224 330500 259000 330528
rect 258224 330488 258230 330500
rect 258994 330488 259000 330500
rect 259052 330488 259058 330540
rect 262398 330488 262404 330540
rect 262456 330528 262462 330540
rect 262582 330528 262588 330540
rect 262456 330500 262588 330528
rect 262456 330488 262462 330500
rect 262582 330488 262588 330500
rect 262640 330488 262646 330540
rect 265158 330488 265164 330540
rect 265216 330528 265222 330540
rect 265894 330528 265900 330540
rect 265216 330500 265900 330528
rect 265216 330488 265222 330500
rect 265894 330488 265900 330500
rect 265952 330488 265958 330540
rect 266446 330488 266452 330540
rect 266504 330528 266510 330540
rect 266998 330528 267004 330540
rect 266504 330500 267004 330528
rect 266504 330488 266510 330500
rect 266998 330488 267004 330500
rect 267056 330488 267062 330540
rect 270586 330488 270592 330540
rect 270644 330528 270650 330540
rect 271322 330528 271328 330540
rect 270644 330500 271328 330528
rect 270644 330488 270650 330500
rect 271322 330488 271328 330500
rect 271380 330488 271386 330540
rect 285766 330488 285772 330540
rect 285824 330528 285830 330540
rect 286318 330528 286324 330540
rect 285824 330500 286324 330528
rect 285824 330488 285830 330500
rect 286318 330488 286324 330500
rect 286376 330488 286382 330540
rect 287146 330488 287152 330540
rect 287204 330528 287210 330540
rect 288158 330528 288164 330540
rect 287204 330500 288164 330528
rect 287204 330488 287210 330500
rect 288158 330488 288164 330500
rect 288216 330488 288222 330540
rect 291286 330488 291292 330540
rect 291344 330528 291350 330540
rect 291838 330528 291844 330540
rect 291344 330500 291844 330528
rect 291344 330488 291350 330500
rect 291838 330488 291844 330500
rect 291896 330488 291902 330540
rect 294046 330488 294052 330540
rect 294104 330528 294110 330540
rect 295150 330528 295156 330540
rect 294104 330500 295156 330528
rect 294104 330488 294110 330500
rect 295150 330488 295156 330500
rect 295208 330488 295214 330540
rect 300946 330488 300952 330540
rect 301004 330528 301010 330540
rect 301682 330528 301688 330540
rect 301004 330500 301688 330528
rect 301004 330488 301010 330500
rect 301682 330488 301688 330500
rect 301740 330488 301746 330540
rect 305086 330488 305092 330540
rect 305144 330528 305150 330540
rect 305730 330528 305736 330540
rect 305144 330500 305736 330528
rect 305144 330488 305150 330500
rect 305730 330488 305736 330500
rect 305788 330488 305794 330540
rect 307754 330488 307760 330540
rect 307812 330528 307818 330540
rect 308582 330528 308588 330540
rect 307812 330500 308588 330528
rect 307812 330488 307818 330500
rect 308582 330488 308588 330500
rect 308640 330488 308646 330540
rect 309318 330488 309324 330540
rect 309376 330528 309382 330540
rect 310054 330528 310060 330540
rect 309376 330500 310060 330528
rect 309376 330488 309382 330500
rect 310054 330488 310060 330500
rect 310112 330488 310118 330540
rect 310606 330488 310612 330540
rect 310664 330528 310670 330540
rect 311158 330528 311164 330540
rect 310664 330500 311164 330528
rect 310664 330488 310670 330500
rect 311158 330488 311164 330500
rect 311216 330488 311222 330540
rect 311986 330488 311992 330540
rect 312044 330528 312050 330540
rect 312630 330528 312636 330540
rect 312044 330500 312636 330528
rect 312044 330488 312050 330500
rect 312630 330488 312636 330500
rect 312688 330488 312694 330540
rect 313274 330488 313280 330540
rect 313332 330528 313338 330540
rect 314102 330528 314108 330540
rect 313332 330500 314108 330528
rect 313332 330488 313338 330500
rect 314102 330488 314108 330500
rect 314160 330488 314166 330540
rect 317598 330488 317604 330540
rect 317656 330528 317662 330540
rect 318518 330528 318524 330540
rect 317656 330500 318524 330528
rect 317656 330488 317662 330500
rect 318518 330488 318524 330500
rect 318576 330488 318582 330540
rect 318886 330488 318892 330540
rect 318944 330528 318950 330540
rect 319530 330528 319536 330540
rect 318944 330500 319536 330528
rect 318944 330488 318950 330500
rect 319530 330488 319536 330500
rect 319588 330488 319594 330540
rect 320266 330488 320272 330540
rect 320324 330528 320330 330540
rect 321002 330528 321008 330540
rect 320324 330500 321008 330528
rect 320324 330488 320330 330500
rect 321002 330488 321008 330500
rect 321060 330488 321066 330540
rect 321646 330488 321652 330540
rect 321704 330528 321710 330540
rect 322106 330528 322112 330540
rect 321704 330500 322112 330528
rect 321704 330488 321710 330500
rect 322106 330488 322112 330500
rect 322164 330488 322170 330540
rect 323118 330488 323124 330540
rect 323176 330528 323182 330540
rect 323946 330528 323952 330540
rect 323176 330500 323952 330528
rect 323176 330488 323182 330500
rect 323946 330488 323952 330500
rect 324004 330488 324010 330540
rect 324498 330488 324504 330540
rect 324556 330528 324562 330540
rect 325418 330528 325424 330540
rect 324556 330500 325424 330528
rect 324556 330488 324562 330500
rect 325418 330488 325424 330500
rect 325476 330488 325482 330540
rect 325786 330488 325792 330540
rect 325844 330528 325850 330540
rect 326522 330528 326528 330540
rect 325844 330500 326528 330528
rect 325844 330488 325850 330500
rect 326522 330488 326528 330500
rect 326580 330488 326586 330540
rect 328546 330488 328552 330540
rect 328604 330528 328610 330540
rect 329466 330528 329472 330540
rect 328604 330500 329472 330528
rect 328604 330488 328610 330500
rect 329466 330488 329472 330500
rect 329524 330488 329530 330540
rect 330018 330488 330024 330540
rect 330076 330528 330082 330540
rect 330570 330528 330576 330540
rect 330076 330500 330576 330528
rect 330076 330488 330082 330500
rect 330570 330488 330576 330500
rect 330628 330488 330634 330540
rect 331306 330488 331312 330540
rect 331364 330528 331370 330540
rect 332318 330528 332324 330540
rect 331364 330500 332324 330528
rect 331364 330488 331370 330500
rect 332318 330488 332324 330500
rect 332376 330488 332382 330540
rect 332686 330488 332692 330540
rect 332744 330528 332750 330540
rect 333422 330528 333428 330540
rect 332744 330500 333428 330528
rect 332744 330488 332750 330500
rect 333422 330488 333428 330500
rect 333480 330488 333486 330540
rect 334066 330488 334072 330540
rect 334124 330528 334130 330540
rect 334526 330528 334532 330540
rect 334124 330500 334532 330528
rect 334124 330488 334130 330500
rect 334526 330488 334532 330500
rect 334584 330488 334590 330540
rect 335538 330488 335544 330540
rect 335596 330528 335602 330540
rect 336366 330528 336372 330540
rect 335596 330500 336372 330528
rect 335596 330488 335602 330500
rect 336366 330488 336372 330500
rect 336424 330488 336430 330540
rect 338114 330488 338120 330540
rect 338172 330528 338178 330540
rect 338942 330528 338948 330540
rect 338172 330500 338948 330528
rect 338172 330488 338178 330500
rect 338942 330488 338948 330500
rect 339000 330488 339006 330540
rect 349982 330488 349988 330540
rect 350040 330528 350046 330540
rect 350442 330528 350448 330540
rect 350040 330500 350448 330528
rect 350040 330488 350046 330500
rect 350442 330488 350448 330500
rect 350500 330488 350506 330540
rect 401870 330488 401876 330540
rect 401928 330528 401934 330540
rect 402790 330528 402796 330540
rect 401928 330500 402796 330528
rect 401928 330488 401934 330500
rect 402790 330488 402796 330500
rect 402848 330488 402854 330540
rect 517514 330528 517520 330540
rect 402946 330500 517520 330528
rect 245654 330460 245660 330472
rect 238726 330432 245660 330460
rect 245654 330420 245660 330432
rect 245712 330420 245718 330472
rect 254026 330420 254032 330472
rect 254084 330460 254090 330472
rect 254946 330460 254952 330472
rect 254084 330432 254952 330460
rect 254084 330420 254090 330432
rect 254946 330420 254952 330432
rect 255004 330420 255010 330472
rect 262306 330420 262312 330472
rect 262364 330460 262370 330472
rect 263318 330460 263324 330472
rect 262364 330432 263324 330460
rect 262364 330420 262370 330432
rect 263318 330420 263324 330432
rect 263376 330420 263382 330472
rect 305178 330420 305184 330472
rect 305236 330460 305242 330472
rect 306098 330460 306104 330472
rect 305236 330432 306104 330460
rect 305236 330420 305242 330432
rect 306098 330420 306104 330432
rect 306156 330420 306162 330472
rect 309134 330420 309140 330472
rect 309192 330460 309198 330472
rect 309686 330460 309692 330472
rect 309192 330432 309692 330460
rect 309192 330420 309198 330432
rect 309686 330420 309692 330432
rect 309744 330420 309750 330472
rect 329926 330420 329932 330472
rect 329984 330460 329990 330472
rect 330938 330460 330944 330472
rect 329984 330432 330944 330460
rect 329984 330420 329990 330432
rect 330938 330420 330944 330432
rect 330996 330420 331002 330472
rect 395246 330420 395252 330472
rect 395304 330460 395310 330472
rect 402946 330460 402974 330500
rect 517514 330488 517520 330500
rect 517572 330488 517578 330540
rect 395304 330432 402974 330460
rect 395304 330420 395310 330432
rect 403250 330420 403256 330472
rect 403308 330460 403314 330472
rect 404170 330460 404176 330472
rect 403308 330432 404176 330460
rect 403308 330420 403314 330432
rect 404170 330420 404176 330432
rect 404228 330420 404234 330472
rect 404722 330420 404728 330472
rect 404780 330460 404786 330472
rect 405458 330460 405464 330472
rect 404780 330432 405464 330460
rect 404780 330420 404786 330432
rect 405458 330420 405464 330432
rect 405516 330420 405522 330472
rect 406194 330420 406200 330472
rect 406252 330460 406258 330472
rect 406930 330460 406936 330472
rect 406252 330432 406936 330460
rect 406252 330420 406258 330432
rect 406930 330420 406936 330432
rect 406988 330420 406994 330472
rect 408770 330420 408776 330472
rect 408828 330460 408834 330472
rect 409690 330460 409696 330472
rect 408828 330432 409696 330460
rect 408828 330420 408834 330432
rect 409690 330420 409696 330432
rect 409748 330420 409754 330472
rect 410242 330420 410248 330472
rect 410300 330460 410306 330472
rect 410978 330460 410984 330472
rect 410300 330432 410984 330460
rect 410300 330420 410306 330432
rect 410978 330420 410984 330432
rect 411036 330420 411042 330472
rect 411714 330420 411720 330472
rect 411772 330460 411778 330472
rect 412542 330460 412548 330472
rect 411772 330432 412548 330460
rect 411772 330420 411778 330432
rect 412542 330420 412548 330432
rect 412600 330420 412606 330472
rect 414290 330420 414296 330472
rect 414348 330460 414354 330472
rect 415210 330460 415216 330472
rect 414348 330432 415216 330460
rect 414348 330420 414354 330432
rect 415210 330420 415216 330432
rect 415268 330420 415274 330472
rect 405090 330352 405096 330404
rect 405148 330392 405154 330404
rect 405642 330392 405648 330404
rect 405148 330364 405648 330392
rect 405148 330352 405154 330364
rect 405642 330352 405648 330364
rect 405700 330352 405706 330404
rect 410610 330352 410616 330404
rect 410668 330392 410674 330404
rect 411162 330392 411168 330404
rect 410668 330364 411168 330392
rect 410668 330352 410674 330364
rect 411162 330352 411168 330364
rect 411220 330352 411226 330404
rect 332594 330148 332600 330200
rect 332652 330188 332658 330200
rect 333054 330188 333060 330200
rect 332652 330160 333060 330188
rect 332652 330148 332658 330160
rect 333054 330148 333060 330160
rect 333112 330148 333118 330200
rect 299566 330012 299572 330064
rect 299624 330052 299630 330064
rect 300578 330052 300584 330064
rect 299624 330024 300584 330052
rect 299624 330012 299630 330024
rect 300578 330012 300584 330024
rect 300636 330012 300642 330064
rect 271966 329808 271972 329860
rect 272024 329848 272030 329860
rect 272426 329848 272432 329860
rect 272024 329820 272432 329848
rect 272024 329808 272030 329820
rect 272426 329808 272432 329820
rect 272484 329808 272490 329860
rect 255314 329604 255320 329656
rect 255372 329644 255378 329656
rect 255682 329644 255688 329656
rect 255372 329616 255688 329644
rect 255372 329604 255378 329616
rect 255682 329604 255688 329616
rect 255740 329604 255746 329656
rect 124122 329400 124128 329452
rect 124180 329440 124186 329452
rect 267734 329440 267740 329452
rect 124180 329412 267740 329440
rect 124180 329400 124186 329412
rect 267734 329400 267740 329412
rect 267792 329400 267798 329452
rect 119982 329332 119988 329384
rect 120040 329372 120046 329384
rect 270034 329372 270040 329384
rect 120040 329344 270040 329372
rect 120040 329332 120046 329344
rect 270034 329332 270040 329344
rect 270092 329332 270098 329384
rect 113082 329264 113088 329316
rect 113140 329304 113146 329316
rect 269574 329304 269580 329316
rect 113140 329276 269580 329304
rect 113140 329264 113146 329276
rect 269574 329264 269580 329276
rect 269632 329264 269638 329316
rect 61378 329196 61384 329248
rect 61436 329236 61442 329248
rect 252554 329236 252560 329248
rect 61436 329208 252560 329236
rect 61436 329196 61442 329208
rect 252554 329196 252560 329208
rect 252612 329196 252618 329248
rect 47578 329128 47584 329180
rect 47636 329168 47642 329180
rect 246574 329168 246580 329180
rect 47636 329140 246580 329168
rect 47636 329128 47642 329140
rect 246574 329128 246580 329140
rect 246632 329128 246638 329180
rect 397362 329128 397368 329180
rect 397420 329168 397426 329180
rect 524414 329168 524420 329180
rect 397420 329140 524420 329168
rect 397420 329128 397426 329140
rect 524414 329128 524420 329140
rect 524472 329128 524478 329180
rect 32398 329060 32404 329112
rect 32456 329100 32462 329112
rect 240318 329100 240324 329112
rect 32456 329072 240324 329100
rect 32456 329060 32462 329072
rect 240318 329060 240324 329072
rect 240376 329060 240382 329112
rect 400766 329060 400772 329112
rect 400824 329100 400830 329112
rect 535454 329100 535460 329112
rect 400824 329072 535460 329100
rect 400824 329060 400830 329072
rect 535454 329060 535460 329072
rect 535512 329060 535518 329112
rect 14458 327700 14464 327752
rect 14516 327740 14522 327752
rect 237742 327740 237748 327752
rect 14516 327712 237748 327740
rect 14516 327700 14522 327712
rect 237742 327700 237748 327712
rect 237800 327700 237806 327752
rect 314746 327156 314752 327208
rect 314804 327196 314810 327208
rect 315574 327196 315580 327208
rect 314804 327168 315580 327196
rect 314804 327156 314810 327168
rect 315574 327156 315580 327168
rect 315632 327156 315638 327208
rect 304994 326884 305000 326936
rect 305052 326924 305058 326936
rect 305362 326924 305368 326936
rect 305052 326896 305368 326924
rect 305052 326884 305058 326896
rect 305362 326884 305368 326896
rect 305420 326884 305426 326936
rect 334158 326680 334164 326732
rect 334216 326720 334222 326732
rect 334894 326720 334900 326732
rect 334216 326692 334900 326720
rect 334216 326680 334222 326692
rect 334894 326680 334900 326692
rect 334952 326680 334958 326732
rect 306466 326476 306472 326528
rect 306524 326516 306530 326528
rect 307478 326516 307484 326528
rect 306524 326488 307484 326516
rect 306524 326476 306530 326488
rect 307478 326476 307484 326488
rect 307536 326476 307542 326528
rect 276198 326408 276204 326460
rect 276256 326408 276262 326460
rect 274634 326340 274640 326392
rect 274692 326380 274698 326392
rect 275738 326380 275744 326392
rect 274692 326352 275744 326380
rect 274692 326340 274698 326352
rect 275738 326340 275744 326352
rect 275796 326340 275802 326392
rect 276216 326256 276244 326408
rect 277486 326340 277492 326392
rect 277544 326380 277550 326392
rect 277670 326380 277676 326392
rect 277544 326352 277676 326380
rect 277544 326340 277550 326352
rect 277670 326340 277676 326352
rect 277728 326340 277734 326392
rect 280246 326340 280252 326392
rect 280304 326380 280310 326392
rect 280890 326380 280896 326392
rect 280304 326352 280896 326380
rect 280304 326340 280310 326352
rect 280890 326340 280896 326352
rect 280948 326340 280954 326392
rect 360930 326340 360936 326392
rect 360988 326380 360994 326392
rect 361298 326380 361304 326392
rect 360988 326352 361304 326380
rect 360988 326340 360994 326352
rect 361298 326340 361304 326352
rect 361356 326340 361362 326392
rect 362402 326340 362408 326392
rect 362460 326380 362466 326392
rect 362862 326380 362868 326392
rect 362460 326352 362868 326380
rect 362460 326340 362466 326352
rect 362862 326340 362868 326352
rect 362920 326340 362926 326392
rect 276198 326204 276204 326256
rect 276256 326204 276262 326256
rect 428550 325592 428556 325644
rect 428608 325632 428614 325644
rect 579890 325632 579896 325644
rect 428608 325604 579896 325632
rect 428608 325592 428614 325604
rect 579890 325592 579896 325604
rect 579948 325592 579954 325644
rect 277486 325116 277492 325168
rect 277544 325156 277550 325168
rect 278314 325156 278320 325168
rect 277544 325128 278320 325156
rect 277544 325116 277550 325128
rect 278314 325116 278320 325128
rect 278372 325116 278378 325168
rect 276106 323620 276112 323672
rect 276164 323660 276170 323672
rect 276290 323660 276296 323672
rect 276164 323632 276296 323660
rect 276164 323620 276170 323632
rect 276290 323620 276296 323632
rect 276348 323620 276354 323672
rect 566458 313216 566464 313268
rect 566516 313256 566522 313268
rect 580166 313256 580172 313268
rect 566516 313228 580172 313256
rect 566516 313216 566522 313228
rect 580166 313216 580172 313228
rect 580224 313216 580230 313268
rect 421650 273164 421656 273216
rect 421708 273204 421714 273216
rect 580166 273204 580172 273216
rect 421708 273176 580172 273204
rect 421708 273164 421714 273176
rect 580166 273164 580172 273176
rect 580224 273164 580230 273216
rect 562318 259360 562324 259412
rect 562376 259400 562382 259412
rect 580166 259400 580172 259412
rect 562376 259372 580172 259400
rect 562376 259360 562382 259372
rect 580166 259360 580172 259372
rect 580224 259360 580230 259412
rect 3326 215228 3332 215280
rect 3384 215268 3390 215280
rect 232590 215268 232596 215280
rect 3384 215240 232596 215268
rect 3384 215228 3390 215240
rect 232590 215228 232596 215240
rect 232648 215228 232654 215280
rect 417418 166948 417424 167000
rect 417476 166988 417482 167000
rect 580166 166988 580172 167000
rect 417476 166960 580172 166988
rect 417476 166948 417482 166960
rect 580166 166948 580172 166960
rect 580224 166948 580230 167000
rect 3418 45500 3424 45552
rect 3476 45540 3482 45552
rect 228358 45540 228364 45552
rect 3476 45512 228364 45540
rect 3476 45500 3482 45512
rect 228358 45500 228364 45512
rect 228416 45500 228422 45552
rect 3418 20612 3424 20664
rect 3476 20652 3482 20664
rect 414934 20652 414940 20664
rect 3476 20624 414940 20652
rect 3476 20612 3482 20624
rect 414934 20612 414940 20624
rect 414992 20612 414998 20664
rect 431218 20612 431224 20664
rect 431276 20652 431282 20664
rect 579982 20652 579988 20664
rect 431276 20624 579988 20652
rect 431276 20612 431282 20624
rect 579982 20612 579988 20624
rect 580040 20612 580046 20664
rect 157242 18572 157248 18624
rect 157300 18612 157306 18624
rect 282178 18612 282184 18624
rect 157300 18584 282184 18612
rect 157300 18572 157306 18584
rect 282178 18572 282184 18584
rect 282236 18572 282242 18624
rect 161290 17212 161296 17264
rect 161348 17252 161354 17264
rect 284386 17252 284392 17264
rect 161348 17224 284392 17252
rect 161348 17212 161354 17224
rect 284386 17212 284392 17224
rect 284444 17212 284450 17264
rect 138842 15852 138848 15904
rect 138900 15892 138906 15904
rect 277578 15892 277584 15904
rect 138900 15864 277584 15892
rect 138900 15852 138906 15864
rect 277578 15852 277584 15864
rect 277636 15852 277642 15904
rect 252370 14424 252376 14476
rect 252428 14464 252434 14476
rect 311986 14464 311992 14476
rect 252428 14436 311992 14464
rect 252428 14424 252434 14436
rect 311986 14424 311992 14436
rect 312044 14424 312050 14476
rect 186130 13336 186136 13388
rect 186188 13376 186194 13388
rect 291286 13376 291292 13388
rect 186188 13348 291292 13376
rect 186188 13336 186194 13348
rect 291286 13336 291292 13348
rect 291344 13336 291350 13388
rect 125870 13268 125876 13320
rect 125928 13308 125934 13320
rect 233970 13308 233976 13320
rect 125928 13280 233976 13308
rect 125928 13268 125934 13280
rect 233970 13268 233976 13280
rect 234028 13268 234034 13320
rect 163682 13200 163688 13252
rect 163740 13240 163746 13252
rect 284478 13240 284484 13252
rect 163740 13212 284484 13240
rect 163740 13200 163746 13212
rect 284478 13200 284484 13212
rect 284536 13200 284542 13252
rect 149514 13132 149520 13184
rect 149572 13172 149578 13184
rect 280246 13172 280252 13184
rect 149572 13144 280252 13172
rect 149572 13132 149578 13144
rect 280246 13132 280252 13144
rect 280304 13132 280310 13184
rect 128170 13064 128176 13116
rect 128228 13104 128234 13116
rect 273438 13104 273444 13116
rect 128228 13076 273444 13104
rect 128228 13064 128234 13076
rect 273438 13064 273444 13076
rect 273496 13064 273502 13116
rect 212166 12180 212172 12232
rect 212224 12220 212230 12232
rect 233878 12220 233884 12232
rect 212224 12192 233884 12220
rect 212224 12180 212230 12192
rect 233878 12180 233884 12192
rect 233936 12180 233942 12232
rect 182542 12112 182548 12164
rect 182600 12152 182606 12164
rect 224218 12152 224224 12164
rect 182600 12124 224224 12152
rect 182600 12112 182606 12124
rect 224218 12112 224224 12124
rect 224276 12112 224282 12164
rect 175458 12044 175464 12096
rect 175516 12084 175522 12096
rect 226978 12084 226984 12096
rect 175516 12056 226984 12084
rect 175516 12044 175522 12056
rect 226978 12044 226984 12056
rect 227036 12044 227042 12096
rect 164878 11976 164884 12028
rect 164936 12016 164942 12028
rect 231118 12016 231124 12028
rect 164936 11988 231124 12016
rect 164936 11976 164942 11988
rect 231118 11976 231124 11988
rect 231176 11976 231182 12028
rect 154206 11908 154212 11960
rect 154264 11948 154270 11960
rect 232498 11948 232504 11960
rect 154264 11920 232504 11948
rect 154264 11908 154270 11920
rect 232498 11908 232504 11920
rect 232556 11908 232562 11960
rect 251082 11908 251088 11960
rect 251140 11948 251146 11960
rect 291838 11948 291844 11960
rect 251140 11920 291844 11948
rect 251140 11908 251146 11920
rect 291838 11908 291844 11920
rect 291896 11908 291902 11960
rect 167178 11840 167184 11892
rect 167236 11880 167242 11892
rect 285766 11880 285772 11892
rect 167236 11852 285772 11880
rect 167236 11840 167242 11852
rect 285766 11840 285772 11852
rect 285824 11840 285830 11892
rect 78582 11772 78588 11824
rect 78640 11812 78646 11824
rect 258350 11812 258356 11824
rect 78640 11784 258356 11812
rect 78640 11772 78646 11784
rect 258350 11772 258356 11784
rect 258408 11772 258414 11824
rect 74442 11704 74448 11756
rect 74500 11744 74506 11756
rect 256878 11744 256884 11756
rect 74500 11716 256884 11744
rect 74500 11704 74506 11716
rect 256878 11704 256884 11716
rect 256936 11704 256942 11756
rect 448606 11704 448612 11756
rect 448664 11744 448670 11756
rect 449802 11744 449808 11756
rect 448664 11716 449808 11744
rect 448664 11704 448670 11716
rect 449802 11704 449808 11716
rect 449860 11704 449866 11756
rect 160094 11636 160100 11688
rect 160152 11676 160158 11688
rect 161290 11676 161296 11688
rect 160152 11648 161296 11676
rect 160152 11636 160158 11648
rect 161290 11636 161296 11648
rect 161348 11636 161354 11688
rect 95050 10956 95056 11008
rect 95108 10996 95114 11008
rect 263686 10996 263692 11008
rect 95108 10968 263692 10996
rect 95108 10956 95114 10968
rect 263686 10956 263692 10968
rect 263744 10956 263750 11008
rect 91002 10888 91008 10940
rect 91060 10928 91066 10940
rect 262398 10928 262404 10940
rect 91060 10900 262404 10928
rect 91060 10888 91066 10900
rect 262398 10888 262404 10900
rect 262456 10888 262462 10940
rect 70302 10820 70308 10872
rect 70360 10860 70366 10872
rect 255590 10860 255596 10872
rect 70360 10832 255596 10860
rect 70360 10820 70366 10832
rect 255590 10820 255596 10832
rect 255648 10820 255654 10872
rect 67542 10752 67548 10804
rect 67600 10792 67606 10804
rect 255498 10792 255504 10804
rect 67600 10764 255504 10792
rect 67600 10752 67606 10764
rect 255498 10752 255504 10764
rect 255556 10752 255562 10804
rect 63218 10684 63224 10736
rect 63276 10724 63282 10736
rect 254210 10724 254216 10736
rect 63276 10696 254216 10724
rect 63276 10684 63282 10696
rect 254210 10684 254216 10696
rect 254268 10684 254274 10736
rect 60642 10616 60648 10668
rect 60700 10656 60706 10668
rect 252738 10656 252744 10668
rect 60700 10628 252744 10656
rect 60700 10616 60706 10628
rect 252738 10616 252744 10628
rect 252796 10616 252802 10668
rect 260650 10616 260656 10668
rect 260708 10656 260714 10668
rect 286318 10656 286324 10668
rect 260708 10628 286324 10656
rect 260708 10616 260714 10628
rect 286318 10616 286324 10628
rect 286376 10616 286382 10668
rect 56502 10548 56508 10600
rect 56560 10588 56566 10600
rect 251266 10588 251272 10600
rect 56560 10560 251272 10588
rect 56560 10548 56566 10560
rect 251266 10548 251272 10560
rect 251324 10548 251330 10600
rect 253474 10548 253480 10600
rect 253532 10588 253538 10600
rect 289078 10588 289084 10600
rect 253532 10560 289084 10588
rect 253532 10548 253538 10560
rect 289078 10548 289084 10560
rect 289136 10548 289142 10600
rect 53742 10480 53748 10532
rect 53800 10520 53806 10532
rect 249886 10520 249892 10532
rect 53800 10492 249892 10520
rect 53800 10480 53806 10492
rect 249886 10480 249892 10492
rect 249944 10480 249950 10532
rect 271782 10480 271788 10532
rect 271840 10520 271846 10532
rect 317598 10520 317604 10532
rect 271840 10492 317604 10520
rect 271840 10480 271846 10492
rect 317598 10480 317604 10492
rect 317656 10480 317662 10532
rect 49602 10412 49608 10464
rect 49660 10452 49666 10464
rect 249978 10452 249984 10464
rect 49660 10424 249984 10452
rect 49660 10412 49666 10424
rect 249978 10412 249984 10424
rect 250036 10412 250042 10464
rect 269022 10412 269028 10464
rect 269080 10452 269086 10464
rect 317506 10452 317512 10464
rect 269080 10424 317512 10452
rect 269080 10412 269086 10424
rect 317506 10412 317512 10424
rect 317564 10412 317570 10464
rect 45462 10344 45468 10396
rect 45520 10384 45526 10396
rect 248598 10384 248604 10396
rect 45520 10356 248604 10384
rect 45520 10344 45526 10356
rect 248598 10344 248604 10356
rect 248656 10344 248662 10396
rect 264882 10344 264888 10396
rect 264940 10384 264946 10396
rect 316126 10384 316132 10396
rect 264940 10356 316132 10384
rect 264940 10344 264946 10356
rect 316126 10344 316132 10356
rect 316184 10344 316190 10396
rect 41322 10276 41328 10328
rect 41380 10316 41386 10328
rect 247126 10316 247132 10328
rect 41380 10288 247132 10316
rect 41380 10276 41386 10288
rect 247126 10276 247132 10288
rect 247184 10276 247190 10328
rect 256602 10276 256608 10328
rect 256660 10316 256666 10328
rect 313458 10316 313464 10328
rect 256660 10288 313464 10316
rect 256660 10276 256666 10288
rect 313458 10276 313464 10288
rect 313516 10276 313522 10328
rect 353018 10276 353024 10328
rect 353076 10316 353082 10328
rect 382366 10316 382372 10328
rect 353076 10288 382372 10316
rect 353076 10276 353082 10288
rect 382366 10276 382372 10288
rect 382424 10276 382430 10328
rect 382918 10276 382924 10328
rect 382976 10316 382982 10328
rect 389450 10316 389456 10328
rect 382976 10288 389456 10316
rect 382976 10276 382982 10288
rect 389450 10276 389456 10288
rect 389508 10276 389514 10328
rect 97902 10208 97908 10260
rect 97960 10248 97966 10260
rect 265066 10248 265072 10260
rect 97960 10220 265072 10248
rect 97960 10208 97966 10220
rect 265066 10208 265072 10220
rect 265124 10208 265130 10260
rect 102042 10140 102048 10192
rect 102100 10180 102106 10192
rect 265158 10180 265164 10192
rect 102100 10152 265164 10180
rect 102100 10140 102106 10152
rect 265158 10140 265164 10152
rect 265216 10140 265222 10192
rect 104526 10072 104532 10124
rect 104584 10112 104590 10124
rect 266446 10112 266452 10124
rect 104584 10084 266452 10112
rect 104584 10072 104590 10084
rect 266446 10072 266452 10084
rect 266504 10072 266510 10124
rect 108942 10004 108948 10056
rect 109000 10044 109006 10056
rect 267826 10044 267832 10056
rect 109000 10016 267832 10044
rect 109000 10004 109006 10016
rect 267826 10004 267832 10016
rect 267884 10004 267890 10056
rect 111610 9936 111616 9988
rect 111668 9976 111674 9988
rect 269298 9976 269304 9988
rect 111668 9948 269304 9976
rect 111668 9936 111674 9948
rect 269298 9936 269304 9948
rect 269356 9936 269362 9988
rect 115842 9868 115848 9920
rect 115900 9908 115906 9920
rect 270678 9908 270684 9920
rect 115900 9880 270684 9908
rect 115900 9868 115906 9880
rect 270678 9868 270684 9880
rect 270736 9868 270742 9920
rect 119798 9800 119804 9852
rect 119856 9840 119862 9852
rect 270586 9840 270592 9852
rect 119856 9812 270592 9840
rect 119856 9800 119862 9812
rect 270586 9800 270592 9812
rect 270644 9800 270650 9852
rect 122742 9732 122748 9784
rect 122800 9772 122806 9784
rect 271966 9772 271972 9784
rect 122800 9744 271972 9772
rect 122800 9732 122806 9744
rect 271966 9732 271972 9744
rect 272024 9732 272030 9784
rect 209774 9596 209780 9648
rect 209832 9636 209838 9648
rect 299658 9636 299664 9648
rect 209832 9608 299664 9636
rect 209832 9596 209838 9608
rect 299658 9596 299664 9608
rect 299716 9596 299722 9648
rect 206186 9528 206192 9580
rect 206244 9568 206250 9580
rect 298186 9568 298192 9580
rect 206244 9540 298192 9568
rect 206244 9528 206250 9540
rect 298186 9528 298192 9540
rect 298244 9528 298250 9580
rect 202690 9460 202696 9512
rect 202748 9500 202754 9512
rect 296806 9500 296812 9512
rect 202748 9472 296812 9500
rect 202748 9460 202754 9472
rect 296806 9460 296812 9472
rect 296864 9460 296870 9512
rect 199102 9392 199108 9444
rect 199160 9432 199166 9444
rect 295518 9432 295524 9444
rect 199160 9404 295524 9432
rect 199160 9392 199166 9404
rect 295518 9392 295524 9404
rect 295576 9392 295582 9444
rect 195606 9324 195612 9376
rect 195664 9364 195670 9376
rect 294046 9364 294052 9376
rect 195664 9336 294052 9364
rect 195664 9324 195670 9336
rect 294046 9324 294052 9336
rect 294104 9324 294110 9376
rect 192018 9256 192024 9308
rect 192076 9296 192082 9308
rect 294138 9296 294144 9308
rect 192076 9268 294144 9296
rect 192076 9256 192082 9268
rect 294138 9256 294144 9268
rect 294196 9256 294202 9308
rect 135254 9188 135260 9240
rect 135312 9228 135318 9240
rect 276106 9228 276112 9240
rect 135312 9200 276112 9228
rect 135312 9188 135318 9200
rect 276106 9188 276112 9200
rect 276164 9188 276170 9240
rect 131758 9120 131764 9172
rect 131816 9160 131822 9172
rect 274910 9160 274916 9172
rect 131816 9132 274916 9160
rect 131816 9120 131822 9132
rect 274910 9120 274916 9132
rect 274968 9120 274974 9172
rect 37182 9052 37188 9104
rect 37240 9092 37246 9104
rect 245838 9092 245844 9104
rect 37240 9064 245844 9092
rect 37240 9052 37246 9064
rect 245838 9052 245844 9064
rect 245896 9052 245902 9104
rect 248782 9052 248788 9104
rect 248840 9092 248846 9104
rect 310790 9092 310796 9104
rect 248840 9064 310796 9092
rect 248840 9052 248846 9064
rect 310790 9052 310796 9064
rect 310848 9052 310854 9104
rect 33594 8984 33600 9036
rect 33652 9024 33658 9036
rect 244366 9024 244372 9036
rect 33652 8996 244372 9024
rect 33652 8984 33658 8996
rect 244366 8984 244372 8996
rect 244424 8984 244430 9036
rect 245194 8984 245200 9036
rect 245252 9024 245258 9036
rect 310698 9024 310704 9036
rect 245252 8996 310704 9024
rect 245252 8984 245258 8996
rect 310698 8984 310704 8996
rect 310756 8984 310762 9036
rect 357158 8984 357164 9036
rect 357216 9024 357222 9036
rect 396534 9024 396540 9036
rect 357216 8996 396540 9024
rect 357216 8984 357222 8996
rect 396534 8984 396540 8996
rect 396592 8984 396598 9036
rect 432598 8984 432604 9036
rect 432656 9024 432662 9036
rect 494698 9024 494704 9036
rect 432656 8996 494704 9024
rect 432656 8984 432662 8996
rect 494698 8984 494704 8996
rect 494756 8984 494762 9036
rect 8754 8916 8760 8968
rect 8812 8956 8818 8968
rect 237466 8956 237472 8968
rect 8812 8928 237472 8956
rect 8812 8916 8818 8928
rect 237466 8916 237472 8928
rect 237524 8916 237530 8968
rect 238110 8916 238116 8968
rect 238168 8956 238174 8968
rect 307938 8956 307944 8968
rect 238168 8928 307944 8956
rect 238168 8916 238174 8928
rect 307938 8916 307944 8928
rect 307996 8916 308002 8968
rect 353938 8916 353944 8968
rect 353996 8956 354002 8968
rect 370590 8956 370596 8968
rect 353996 8928 370596 8956
rect 353996 8916 354002 8928
rect 370590 8916 370596 8928
rect 370648 8916 370654 8968
rect 372430 8916 372436 8968
rect 372488 8956 372494 8968
rect 445018 8956 445024 8968
rect 372488 8928 445024 8956
rect 372488 8916 372494 8928
rect 445018 8916 445024 8928
rect 445076 8916 445082 8968
rect 126974 8848 126980 8900
rect 127032 8888 127038 8900
rect 213178 8888 213184 8900
rect 127032 8860 213184 8888
rect 127032 8848 127038 8860
rect 213178 8848 213184 8860
rect 213236 8848 213242 8900
rect 213362 8848 213368 8900
rect 213420 8888 213426 8900
rect 299566 8888 299572 8900
rect 213420 8860 299572 8888
rect 213420 8848 213426 8860
rect 299566 8848 299572 8860
rect 299624 8848 299630 8900
rect 216858 8780 216864 8832
rect 216916 8820 216922 8832
rect 300946 8820 300952 8832
rect 216916 8792 300952 8820
rect 216916 8780 216922 8792
rect 300946 8780 300952 8792
rect 301004 8780 301010 8832
rect 220446 8712 220452 8764
rect 220504 8752 220510 8764
rect 302418 8752 302424 8764
rect 220504 8724 302424 8752
rect 220504 8712 220510 8724
rect 302418 8712 302424 8724
rect 302476 8712 302482 8764
rect 223942 8644 223948 8696
rect 224000 8684 224006 8696
rect 303706 8684 303712 8696
rect 224000 8656 303712 8684
rect 224000 8644 224006 8656
rect 303706 8644 303712 8656
rect 303764 8644 303770 8696
rect 227530 8576 227536 8628
rect 227588 8616 227594 8628
rect 305270 8616 305276 8628
rect 227588 8588 305276 8616
rect 227588 8576 227594 8588
rect 305270 8576 305276 8588
rect 305328 8576 305334 8628
rect 231026 8508 231032 8560
rect 231084 8548 231090 8560
rect 305178 8548 305184 8560
rect 231084 8520 305184 8548
rect 231084 8508 231090 8520
rect 305178 8508 305184 8520
rect 305236 8508 305242 8560
rect 234982 8440 234988 8492
rect 235040 8480 235046 8492
rect 306650 8480 306656 8492
rect 235040 8452 306656 8480
rect 235040 8440 235046 8452
rect 306650 8440 306656 8452
rect 306708 8440 306714 8492
rect 241698 8372 241704 8424
rect 241756 8412 241762 8424
rect 309410 8412 309416 8424
rect 241756 8384 309416 8412
rect 241756 8372 241762 8384
rect 309410 8372 309416 8384
rect 309468 8372 309474 8424
rect 421558 8304 421564 8356
rect 421616 8344 421622 8356
rect 423766 8344 423772 8356
rect 421616 8316 423772 8344
rect 421616 8304 421622 8316
rect 423766 8304 423772 8316
rect 423824 8304 423830 8356
rect 428458 8304 428464 8356
rect 428516 8344 428522 8356
rect 434438 8344 434444 8356
rect 428516 8316 434444 8344
rect 428516 8304 428522 8316
rect 434438 8304 434444 8316
rect 434496 8304 434502 8356
rect 137646 8236 137652 8288
rect 137704 8276 137710 8288
rect 277670 8276 277676 8288
rect 137704 8248 277676 8276
rect 137704 8236 137710 8248
rect 277670 8236 277676 8248
rect 277728 8236 277734 8288
rect 372338 8236 372344 8288
rect 372396 8276 372402 8288
rect 442626 8276 442632 8288
rect 372396 8248 442632 8276
rect 372396 8236 372402 8248
rect 442626 8236 442632 8248
rect 442684 8236 442690 8288
rect 134150 8168 134156 8220
rect 134208 8208 134214 8220
rect 276198 8208 276204 8220
rect 134208 8180 276204 8208
rect 134208 8168 134214 8180
rect 276198 8168 276204 8180
rect 276256 8168 276262 8220
rect 403986 8168 403992 8220
rect 404044 8208 404050 8220
rect 545482 8208 545488 8220
rect 404044 8180 545488 8208
rect 404044 8168 404050 8180
rect 545482 8168 545488 8180
rect 545540 8168 545546 8220
rect 79686 8100 79692 8152
rect 79744 8140 79750 8152
rect 258077 8143 258135 8149
rect 258077 8140 258089 8143
rect 79744 8112 258089 8140
rect 79744 8100 79750 8112
rect 258077 8109 258089 8112
rect 258123 8109 258135 8143
rect 258350 8140 258356 8152
rect 258077 8103 258135 8109
rect 258184 8112 258356 8140
rect 76190 8032 76196 8084
rect 76248 8072 76254 8084
rect 258184 8072 258212 8112
rect 258350 8100 258356 8112
rect 258408 8100 258414 8152
rect 258445 8143 258503 8149
rect 258445 8109 258457 8143
rect 258491 8140 258503 8143
rect 259546 8140 259552 8152
rect 258491 8112 259552 8140
rect 258491 8109 258503 8112
rect 258445 8103 258503 8109
rect 259546 8100 259552 8112
rect 259604 8100 259610 8152
rect 265342 8100 265348 8152
rect 265400 8140 265406 8152
rect 316218 8140 316224 8152
rect 265400 8112 316224 8140
rect 265400 8100 265406 8112
rect 316218 8100 316224 8112
rect 316276 8100 316282 8152
rect 405458 8100 405464 8152
rect 405516 8140 405522 8152
rect 549070 8140 549076 8152
rect 405516 8112 549076 8140
rect 405516 8100 405522 8112
rect 549070 8100 549076 8112
rect 549128 8100 549134 8152
rect 76248 8044 258212 8072
rect 76248 8032 76254 8044
rect 258258 8032 258264 8084
rect 258316 8072 258322 8084
rect 258316 8044 261064 8072
rect 258316 8032 258322 8044
rect 72602 7964 72608 8016
rect 72660 8004 72666 8016
rect 256786 8004 256792 8016
rect 72660 7976 256792 8004
rect 72660 7964 72666 7976
rect 256786 7964 256792 7976
rect 256844 7964 256850 8016
rect 258077 8007 258135 8013
rect 258077 7973 258089 8007
rect 258123 8004 258135 8007
rect 261036 8004 261064 8044
rect 261754 8032 261760 8084
rect 261812 8072 261818 8084
rect 314746 8072 314752 8084
rect 261812 8044 314752 8072
rect 261812 8032 261818 8044
rect 314746 8032 314752 8044
rect 314804 8032 314810 8084
rect 405366 8032 405372 8084
rect 405424 8072 405430 8084
rect 552658 8072 552664 8084
rect 405424 8044 552664 8072
rect 405424 8032 405430 8044
rect 552658 8032 552664 8044
rect 552716 8032 552722 8084
rect 314838 8004 314844 8016
rect 258123 7976 258304 8004
rect 261036 7976 314844 8004
rect 258123 7973 258135 7976
rect 258077 7967 258135 7973
rect 30098 7896 30104 7948
rect 30156 7936 30162 7948
rect 243078 7936 243084 7948
rect 30156 7908 243084 7936
rect 30156 7896 30162 7908
rect 243078 7896 243084 7908
rect 243136 7896 243142 7948
rect 251174 7896 251180 7948
rect 251232 7936 251238 7948
rect 258276 7936 258304 7976
rect 314838 7964 314844 7976
rect 314896 7964 314902 8016
rect 406746 7964 406752 8016
rect 406804 8004 406810 8016
rect 556154 8004 556160 8016
rect 406804 7976 556160 8004
rect 406804 7964 406810 7976
rect 556154 7964 556160 7976
rect 556212 7964 556218 8016
rect 313366 7936 313372 7948
rect 251232 7908 258212 7936
rect 258276 7908 313372 7936
rect 251232 7896 251238 7908
rect 26510 7828 26516 7880
rect 26568 7868 26574 7880
rect 242986 7868 242992 7880
rect 26568 7840 242992 7868
rect 26568 7828 26574 7840
rect 242986 7828 242992 7840
rect 243044 7828 243050 7880
rect 254670 7828 254676 7880
rect 254728 7868 254734 7880
rect 258077 7871 258135 7877
rect 258077 7868 258089 7871
rect 254728 7840 258089 7868
rect 254728 7828 254734 7840
rect 258077 7837 258089 7840
rect 258123 7837 258135 7871
rect 258184 7868 258212 7908
rect 313366 7896 313372 7908
rect 313424 7896 313430 7948
rect 408218 7896 408224 7948
rect 408276 7936 408282 7948
rect 559742 7936 559748 7948
rect 408276 7908 559748 7936
rect 408276 7896 408282 7908
rect 559742 7896 559748 7908
rect 559800 7896 559806 7948
rect 312078 7868 312084 7880
rect 258184 7840 312084 7868
rect 258077 7831 258135 7837
rect 312078 7828 312084 7840
rect 312136 7828 312142 7880
rect 409506 7828 409512 7880
rect 409564 7868 409570 7880
rect 563238 7868 563244 7880
rect 409564 7840 563244 7868
rect 409564 7828 409570 7840
rect 563238 7828 563244 7840
rect 563296 7828 563302 7880
rect 21818 7760 21824 7812
rect 21876 7800 21882 7812
rect 241790 7800 241796 7812
rect 21876 7772 241796 7800
rect 21876 7760 21882 7772
rect 241790 7760 241796 7772
rect 241848 7760 241854 7812
rect 247586 7760 247592 7812
rect 247644 7800 247650 7812
rect 310606 7800 310612 7812
rect 247644 7772 310612 7800
rect 247644 7760 247650 7772
rect 310606 7760 310612 7772
rect 310664 7760 310670 7812
rect 410978 7760 410984 7812
rect 411036 7800 411042 7812
rect 566826 7800 566832 7812
rect 411036 7772 566832 7800
rect 411036 7760 411042 7772
rect 566826 7760 566832 7772
rect 566884 7760 566890 7812
rect 17034 7692 17040 7744
rect 17092 7732 17098 7744
rect 240134 7732 240140 7744
rect 17092 7704 240140 7732
rect 17092 7692 17098 7704
rect 240134 7692 240140 7704
rect 240192 7692 240198 7744
rect 244090 7692 244096 7744
rect 244148 7732 244154 7744
rect 309318 7732 309324 7744
rect 244148 7704 309324 7732
rect 244148 7692 244154 7704
rect 309318 7692 309324 7704
rect 309376 7692 309382 7744
rect 410886 7692 410892 7744
rect 410944 7732 410950 7744
rect 570322 7732 570328 7744
rect 410944 7704 570328 7732
rect 410944 7692 410950 7704
rect 570322 7692 570328 7704
rect 570380 7692 570386 7744
rect 12342 7624 12348 7676
rect 12400 7664 12406 7676
rect 237374 7664 237380 7676
rect 12400 7636 237380 7664
rect 12400 7624 12406 7636
rect 237374 7624 237380 7636
rect 237432 7624 237438 7676
rect 240502 7624 240508 7676
rect 240560 7664 240566 7676
rect 309226 7664 309232 7676
rect 240560 7636 309232 7664
rect 240560 7624 240566 7636
rect 309226 7624 309232 7636
rect 309284 7624 309290 7676
rect 412266 7624 412272 7676
rect 412324 7664 412330 7676
rect 573910 7664 573916 7676
rect 412324 7636 573916 7664
rect 412324 7624 412330 7636
rect 573910 7624 573916 7636
rect 573968 7624 573974 7676
rect 4062 7556 4068 7608
rect 4120 7596 4126 7608
rect 236178 7596 236184 7608
rect 4120 7568 236184 7596
rect 4120 7556 4126 7568
rect 236178 7556 236184 7568
rect 236236 7556 236242 7608
rect 237006 7556 237012 7608
rect 237064 7596 237070 7608
rect 307846 7596 307852 7608
rect 237064 7568 307852 7596
rect 237064 7556 237070 7568
rect 307846 7556 307852 7568
rect 307904 7556 307910 7608
rect 413738 7556 413744 7608
rect 413796 7596 413802 7608
rect 577406 7596 577412 7608
rect 413796 7568 577412 7596
rect 413796 7556 413802 7568
rect 577406 7556 577412 7568
rect 577464 7556 577470 7608
rect 141234 7488 141240 7540
rect 141292 7528 141298 7540
rect 277486 7528 277492 7540
rect 141292 7500 277492 7528
rect 141292 7488 141298 7500
rect 277486 7488 277492 7500
rect 277544 7488 277550 7540
rect 371050 7488 371056 7540
rect 371108 7528 371114 7540
rect 371108 7500 435312 7528
rect 371108 7488 371114 7500
rect 144730 7420 144736 7472
rect 144788 7460 144794 7472
rect 278958 7460 278964 7472
rect 144788 7432 278964 7460
rect 144788 7420 144794 7432
rect 278958 7420 278964 7432
rect 279016 7420 279022 7472
rect 369670 7420 369676 7472
rect 369728 7460 369734 7472
rect 369728 7432 433748 7460
rect 369728 7420 369734 7432
rect 148318 7352 148324 7404
rect 148376 7392 148382 7404
rect 280338 7392 280344 7404
rect 148376 7364 280344 7392
rect 148376 7352 148382 7364
rect 280338 7352 280344 7364
rect 280396 7352 280402 7404
rect 368198 7352 368204 7404
rect 368256 7392 368262 7404
rect 432046 7392 432052 7404
rect 368256 7364 432052 7392
rect 368256 7352 368262 7364
rect 432046 7352 432052 7364
rect 432104 7352 432110 7404
rect 151814 7284 151820 7336
rect 151872 7324 151878 7336
rect 281718 7324 281724 7336
rect 151872 7296 281724 7324
rect 151872 7284 151878 7296
rect 281718 7284 281724 7296
rect 281776 7284 281782 7336
rect 368290 7284 368296 7336
rect 368348 7324 368354 7336
rect 368348 7296 425376 7324
rect 368348 7284 368354 7296
rect 155402 7216 155408 7268
rect 155460 7256 155466 7268
rect 283006 7256 283012 7268
rect 155460 7228 283012 7256
rect 155460 7216 155466 7228
rect 283006 7216 283012 7228
rect 283064 7216 283070 7268
rect 367002 7216 367008 7268
rect 367060 7256 367066 7268
rect 424962 7256 424968 7268
rect 367060 7228 424968 7256
rect 367060 7216 367066 7228
rect 424962 7216 424968 7228
rect 425020 7216 425026 7268
rect 425348 7256 425376 7296
rect 425698 7284 425704 7336
rect 425756 7324 425762 7336
rect 427262 7324 427268 7336
rect 425756 7296 427268 7324
rect 425756 7284 425762 7296
rect 427262 7284 427268 7296
rect 427320 7284 427326 7336
rect 433720 7324 433748 7432
rect 435284 7392 435312 7500
rect 435358 7488 435364 7540
rect 435416 7528 435422 7540
rect 437934 7528 437940 7540
rect 435416 7500 437940 7528
rect 435416 7488 435422 7500
rect 437934 7488 437940 7500
rect 437992 7488 437998 7540
rect 439130 7392 439136 7404
rect 435284 7364 439136 7392
rect 439130 7352 439136 7364
rect 439188 7352 439194 7404
rect 435542 7324 435548 7336
rect 433720 7296 435548 7324
rect 435542 7284 435548 7296
rect 435600 7284 435606 7336
rect 428458 7256 428464 7268
rect 425348 7228 428464 7256
rect 428458 7216 428464 7228
rect 428516 7216 428522 7268
rect 158898 7148 158904 7200
rect 158956 7188 158962 7200
rect 283098 7188 283104 7200
rect 158956 7160 283104 7188
rect 158956 7148 158962 7160
rect 283098 7148 283104 7160
rect 283156 7148 283162 7200
rect 365530 7148 365536 7200
rect 365588 7188 365594 7200
rect 421374 7188 421380 7200
rect 365588 7160 421380 7188
rect 365588 7148 365594 7160
rect 421374 7148 421380 7160
rect 421432 7148 421438 7200
rect 229830 7080 229836 7132
rect 229888 7120 229894 7132
rect 305086 7120 305092 7132
rect 229888 7092 305092 7120
rect 229888 7080 229894 7092
rect 305086 7080 305092 7092
rect 305144 7080 305150 7132
rect 364150 7080 364156 7132
rect 364208 7120 364214 7132
rect 417878 7120 417884 7132
rect 364208 7092 417884 7120
rect 364208 7080 364214 7092
rect 417878 7080 417884 7092
rect 417936 7080 417942 7132
rect 233418 7012 233424 7064
rect 233476 7052 233482 7064
rect 306558 7052 306564 7064
rect 233476 7024 306564 7052
rect 233476 7012 233482 7024
rect 306558 7012 306564 7024
rect 306616 7012 306622 7064
rect 362586 7012 362592 7064
rect 362644 7052 362650 7064
rect 414290 7052 414296 7064
rect 362644 7024 414296 7052
rect 362644 7012 362650 7024
rect 414290 7012 414296 7024
rect 414348 7012 414354 7064
rect 234614 6808 234620 6860
rect 234672 6848 234678 6860
rect 580166 6848 580172 6860
rect 234672 6820 580172 6848
rect 234672 6808 234678 6820
rect 580166 6808 580172 6820
rect 580224 6808 580230 6860
rect 169570 6740 169576 6792
rect 169628 6780 169634 6792
rect 287238 6780 287244 6792
rect 169628 6752 287244 6780
rect 169628 6740 169634 6752
rect 287238 6740 287244 6752
rect 287296 6740 287302 6792
rect 382090 6740 382096 6792
rect 382148 6780 382154 6792
rect 476942 6780 476948 6792
rect 382148 6752 476948 6780
rect 382148 6740 382154 6752
rect 476942 6740 476948 6752
rect 477000 6740 477006 6792
rect 166074 6672 166080 6724
rect 166132 6712 166138 6724
rect 285858 6712 285864 6724
rect 166132 6684 285864 6712
rect 166132 6672 166138 6684
rect 285858 6672 285864 6684
rect 285916 6672 285922 6724
rect 384850 6672 384856 6724
rect 384908 6712 384914 6724
rect 481726 6712 481732 6724
rect 384908 6684 481732 6712
rect 384908 6672 384914 6684
rect 481726 6672 481732 6684
rect 481784 6672 481790 6724
rect 130562 6604 130568 6656
rect 130620 6644 130626 6656
rect 274818 6644 274824 6656
rect 130620 6616 274824 6644
rect 130620 6604 130626 6616
rect 274818 6604 274824 6616
rect 274876 6604 274882 6656
rect 384758 6604 384764 6656
rect 384816 6644 384822 6656
rect 485222 6644 485228 6656
rect 384816 6616 485228 6644
rect 384816 6604 384822 6616
rect 485222 6604 485228 6616
rect 485280 6604 485286 6656
rect 69106 6536 69112 6588
rect 69164 6576 69170 6588
rect 255406 6576 255412 6588
rect 69164 6548 255412 6576
rect 69164 6536 69170 6548
rect 255406 6536 255412 6548
rect 255464 6536 255470 6588
rect 386322 6536 386328 6588
rect 386380 6576 386386 6588
rect 488810 6576 488816 6588
rect 386380 6548 488816 6576
rect 386380 6536 386386 6548
rect 488810 6536 488816 6548
rect 488868 6536 488874 6588
rect 65518 6468 65524 6520
rect 65576 6508 65582 6520
rect 254026 6508 254032 6520
rect 65576 6480 254032 6508
rect 65576 6468 65582 6480
rect 254026 6468 254032 6480
rect 254084 6468 254090 6520
rect 387702 6468 387708 6520
rect 387760 6508 387766 6520
rect 492306 6508 492312 6520
rect 387760 6480 492312 6508
rect 387760 6468 387766 6480
rect 492306 6468 492312 6480
rect 492364 6468 492370 6520
rect 62022 6400 62028 6452
rect 62080 6440 62086 6452
rect 254118 6440 254124 6452
rect 62080 6412 254124 6440
rect 62080 6400 62086 6412
rect 254118 6400 254124 6412
rect 254176 6400 254182 6452
rect 389082 6400 389088 6452
rect 389140 6440 389146 6452
rect 495894 6440 495900 6452
rect 389140 6412 495900 6440
rect 389140 6400 389146 6412
rect 495894 6400 495900 6412
rect 495952 6400 495958 6452
rect 58434 6332 58440 6384
rect 58492 6372 58498 6384
rect 252646 6372 252652 6384
rect 58492 6344 252652 6372
rect 58492 6332 58498 6344
rect 252646 6332 252652 6344
rect 252704 6332 252710 6384
rect 299658 6332 299664 6384
rect 299716 6372 299722 6384
rect 316678 6372 316684 6384
rect 299716 6344 316684 6372
rect 299716 6332 299722 6344
rect 316678 6332 316684 6344
rect 316736 6332 316742 6384
rect 390186 6332 390192 6384
rect 390244 6372 390250 6384
rect 499390 6372 499396 6384
rect 390244 6344 499396 6372
rect 390244 6332 390250 6344
rect 499390 6332 499396 6344
rect 499448 6332 499454 6384
rect 54938 6264 54944 6316
rect 54996 6304 55002 6316
rect 251358 6304 251364 6316
rect 54996 6276 251364 6304
rect 54996 6264 55002 6276
rect 251358 6264 251364 6276
rect 251416 6264 251422 6316
rect 259454 6264 259460 6316
rect 259512 6304 259518 6316
rect 295978 6304 295984 6316
rect 259512 6276 295984 6304
rect 259512 6264 259518 6276
rect 295978 6264 295984 6276
rect 296036 6264 296042 6316
rect 303154 6264 303160 6316
rect 303212 6304 303218 6316
rect 327718 6304 327724 6316
rect 303212 6276 327724 6304
rect 303212 6264 303218 6276
rect 327718 6264 327724 6276
rect 327776 6264 327782 6316
rect 390370 6264 390376 6316
rect 390428 6304 390434 6316
rect 502886 6304 502892 6316
rect 390428 6276 502892 6304
rect 390428 6264 390434 6276
rect 502886 6264 502892 6276
rect 502944 6264 502950 6316
rect 51350 6196 51356 6248
rect 51408 6236 51414 6248
rect 250070 6236 250076 6248
rect 51408 6208 250076 6236
rect 51408 6196 51414 6208
rect 250070 6196 250076 6208
rect 250128 6196 250134 6248
rect 268838 6196 268844 6248
rect 268896 6236 268902 6248
rect 317690 6236 317696 6248
rect 268896 6208 317696 6236
rect 268896 6196 268902 6208
rect 317690 6196 317696 6208
rect 317748 6196 317754 6248
rect 371878 6196 371884 6248
rect 371936 6236 371942 6248
rect 378870 6236 378876 6248
rect 371936 6208 378876 6236
rect 371936 6196 371942 6208
rect 378870 6196 378876 6208
rect 378928 6196 378934 6248
rect 391658 6196 391664 6248
rect 391716 6236 391722 6248
rect 506566 6236 506572 6248
rect 391716 6208 506572 6236
rect 391716 6196 391722 6208
rect 506566 6196 506572 6208
rect 506624 6196 506630 6248
rect 47854 6128 47860 6180
rect 47912 6168 47918 6180
rect 248506 6168 248512 6180
rect 47912 6140 248512 6168
rect 47912 6128 47918 6140
rect 248506 6128 248512 6140
rect 248564 6128 248570 6180
rect 257062 6128 257068 6180
rect 257120 6168 257126 6180
rect 313274 6168 313280 6180
rect 257120 6140 313280 6168
rect 257120 6128 257126 6140
rect 313274 6128 313280 6140
rect 313332 6128 313338 6180
rect 370498 6128 370504 6180
rect 370556 6168 370562 6180
rect 385954 6168 385960 6180
rect 370556 6140 385960 6168
rect 370556 6128 370562 6140
rect 385954 6128 385960 6140
rect 386012 6128 386018 6180
rect 393130 6128 393136 6180
rect 393188 6168 393194 6180
rect 510062 6168 510068 6180
rect 393188 6140 510068 6168
rect 393188 6128 393194 6140
rect 510062 6128 510068 6140
rect 510120 6128 510126 6180
rect 173158 6060 173164 6112
rect 173216 6100 173222 6112
rect 287146 6100 287152 6112
rect 173216 6072 287152 6100
rect 173216 6060 173222 6072
rect 287146 6060 287152 6072
rect 287204 6060 287210 6112
rect 381998 6060 382004 6112
rect 382056 6100 382062 6112
rect 473446 6100 473452 6112
rect 382056 6072 473452 6100
rect 382056 6060 382062 6072
rect 473446 6060 473452 6072
rect 473504 6060 473510 6112
rect 176654 5992 176660 6044
rect 176712 6032 176718 6044
rect 288618 6032 288624 6044
rect 176712 6004 288624 6032
rect 176712 5992 176718 6004
rect 288618 5992 288624 6004
rect 288676 5992 288682 6044
rect 380710 5992 380716 6044
rect 380768 6032 380774 6044
rect 469858 6032 469864 6044
rect 380768 6004 469864 6032
rect 380768 5992 380774 6004
rect 469858 5992 469864 6004
rect 469916 5992 469922 6044
rect 180242 5924 180248 5976
rect 180300 5964 180306 5976
rect 289998 5964 290004 5976
rect 180300 5936 290004 5964
rect 180300 5924 180306 5936
rect 289998 5924 290004 5936
rect 290056 5924 290062 5976
rect 379422 5924 379428 5976
rect 379480 5964 379486 5976
rect 466270 5964 466276 5976
rect 379480 5936 466276 5964
rect 379480 5924 379486 5936
rect 466270 5924 466276 5936
rect 466328 5924 466334 5976
rect 468478 5924 468484 5976
rect 468536 5964 468542 5976
rect 474550 5964 474556 5976
rect 468536 5936 474556 5964
rect 468536 5924 468542 5936
rect 474550 5924 474556 5936
rect 474608 5924 474614 5976
rect 183738 5856 183744 5908
rect 183796 5896 183802 5908
rect 291378 5896 291384 5908
rect 183796 5868 291384 5896
rect 183796 5856 183802 5868
rect 291378 5856 291384 5868
rect 291436 5856 291442 5908
rect 377950 5856 377956 5908
rect 378008 5896 378014 5908
rect 462774 5896 462780 5908
rect 378008 5868 462780 5896
rect 378008 5856 378014 5868
rect 462774 5856 462780 5868
rect 462832 5856 462838 5908
rect 187326 5788 187332 5840
rect 187384 5828 187390 5840
rect 292666 5828 292672 5840
rect 187384 5800 292672 5828
rect 187384 5788 187390 5800
rect 292666 5788 292672 5800
rect 292724 5788 292730 5840
rect 377858 5788 377864 5840
rect 377916 5828 377922 5840
rect 459186 5828 459192 5840
rect 377916 5800 459192 5828
rect 377916 5788 377922 5800
rect 459186 5788 459192 5800
rect 459244 5788 459250 5840
rect 190822 5720 190828 5772
rect 190880 5760 190886 5772
rect 292758 5760 292764 5772
rect 190880 5732 292764 5760
rect 190880 5720 190886 5732
rect 292758 5720 292764 5732
rect 292816 5720 292822 5772
rect 376662 5720 376668 5772
rect 376720 5760 376726 5772
rect 455690 5760 455696 5772
rect 376720 5732 455696 5760
rect 376720 5720 376726 5732
rect 455690 5720 455696 5732
rect 455748 5720 455754 5772
rect 194410 5652 194416 5704
rect 194468 5692 194474 5704
rect 294230 5692 294236 5704
rect 194468 5664 294236 5692
rect 194468 5652 194474 5664
rect 294230 5652 294236 5664
rect 294288 5652 294294 5704
rect 375190 5652 375196 5704
rect 375248 5692 375254 5704
rect 452102 5692 452108 5704
rect 375248 5664 452108 5692
rect 375248 5652 375254 5664
rect 452102 5652 452108 5664
rect 452160 5652 452166 5704
rect 363598 5516 363604 5568
rect 363656 5556 363662 5568
rect 367002 5556 367008 5568
rect 363656 5528 367008 5556
rect 363656 5516 363662 5528
rect 367002 5516 367008 5528
rect 367060 5516 367066 5568
rect 475378 5516 475384 5568
rect 475436 5556 475442 5568
rect 480530 5556 480536 5568
rect 475436 5528 480536 5556
rect 475436 5516 475442 5528
rect 480530 5516 480536 5528
rect 480588 5516 480594 5568
rect 486510 5516 486516 5568
rect 486568 5556 486574 5568
rect 487614 5556 487620 5568
rect 486568 5528 487620 5556
rect 486568 5516 486574 5528
rect 487614 5516 487620 5528
rect 487672 5516 487678 5568
rect 497458 5516 497464 5568
rect 497516 5556 497522 5568
rect 498194 5556 498200 5568
rect 497516 5528 498200 5556
rect 497516 5516 497522 5528
rect 498194 5516 498200 5528
rect 498252 5516 498258 5568
rect 504358 5516 504364 5568
rect 504416 5556 504422 5568
rect 505370 5556 505376 5568
rect 504416 5528 505376 5556
rect 504416 5516 504422 5528
rect 505370 5516 505376 5528
rect 505428 5516 505434 5568
rect 186222 5448 186228 5500
rect 186280 5488 186286 5500
rect 215938 5488 215944 5500
rect 186280 5460 215944 5488
rect 186280 5448 186286 5460
rect 215938 5448 215944 5460
rect 215996 5448 216002 5500
rect 218054 5448 218060 5500
rect 218112 5488 218118 5500
rect 302326 5488 302332 5500
rect 218112 5460 302332 5488
rect 218112 5448 218118 5460
rect 302326 5448 302332 5460
rect 302384 5448 302390 5500
rect 355778 5448 355784 5500
rect 355836 5488 355842 5500
rect 391842 5488 391848 5500
rect 355836 5460 391848 5488
rect 355836 5448 355842 5460
rect 391842 5448 391848 5460
rect 391900 5448 391906 5500
rect 402698 5448 402704 5500
rect 402756 5488 402762 5500
rect 540790 5488 540796 5500
rect 402756 5460 540796 5488
rect 402756 5448 402762 5460
rect 540790 5448 540796 5460
rect 540848 5448 540854 5500
rect 189718 5380 189724 5432
rect 189776 5420 189782 5432
rect 214282 5420 214288 5432
rect 189776 5392 214288 5420
rect 189776 5380 189782 5392
rect 214282 5380 214288 5392
rect 214340 5380 214346 5432
rect 214466 5380 214472 5432
rect 214524 5420 214530 5432
rect 301038 5420 301044 5432
rect 214524 5392 301044 5420
rect 214524 5380 214530 5392
rect 301038 5380 301044 5392
rect 301096 5380 301102 5432
rect 357250 5380 357256 5432
rect 357308 5420 357314 5432
rect 395338 5420 395344 5432
rect 357308 5392 395344 5420
rect 357308 5380 357314 5392
rect 395338 5380 395344 5392
rect 395396 5380 395402 5432
rect 404170 5380 404176 5432
rect 404228 5420 404234 5432
rect 544378 5420 544384 5432
rect 404228 5392 544384 5420
rect 404228 5380 404234 5392
rect 544378 5380 544384 5392
rect 544436 5380 544442 5432
rect 210970 5312 210976 5364
rect 211028 5352 211034 5364
rect 299750 5352 299756 5364
rect 211028 5324 299756 5352
rect 211028 5312 211034 5324
rect 299750 5312 299756 5324
rect 299808 5312 299814 5364
rect 358538 5312 358544 5364
rect 358596 5352 358602 5364
rect 400122 5352 400128 5364
rect 358596 5324 400128 5352
rect 358596 5312 358602 5324
rect 400122 5312 400128 5324
rect 400180 5312 400186 5364
rect 404078 5312 404084 5364
rect 404136 5352 404142 5364
rect 547874 5352 547880 5364
rect 404136 5324 547880 5352
rect 404136 5312 404142 5324
rect 547874 5312 547880 5324
rect 547932 5312 547938 5364
rect 136450 5244 136456 5296
rect 136508 5284 136514 5296
rect 204898 5284 204904 5296
rect 136508 5256 204904 5284
rect 136508 5244 136514 5256
rect 204898 5244 204904 5256
rect 204956 5244 204962 5296
rect 207382 5244 207388 5296
rect 207440 5284 207446 5296
rect 298278 5284 298284 5296
rect 207440 5256 298284 5284
rect 207440 5244 207446 5256
rect 298278 5244 298284 5256
rect 298336 5244 298342 5296
rect 358630 5244 358636 5296
rect 358688 5284 358694 5296
rect 398926 5284 398932 5296
rect 358688 5256 398932 5284
rect 358688 5244 358694 5256
rect 398926 5244 398932 5256
rect 398984 5244 398990 5296
rect 405550 5244 405556 5296
rect 405608 5284 405614 5296
rect 551462 5284 551468 5296
rect 405608 5256 551468 5284
rect 405608 5244 405614 5256
rect 551462 5244 551468 5256
rect 551520 5244 551526 5296
rect 203886 5176 203892 5228
rect 203944 5216 203950 5228
rect 296898 5216 296904 5228
rect 203944 5188 296904 5216
rect 203944 5176 203950 5188
rect 296898 5176 296904 5188
rect 296956 5176 296962 5228
rect 359826 5176 359832 5228
rect 359884 5216 359890 5228
rect 402514 5216 402520 5228
rect 359884 5188 402520 5216
rect 359884 5176 359890 5188
rect 402514 5176 402520 5188
rect 402572 5176 402578 5228
rect 406838 5176 406844 5228
rect 406896 5216 406902 5228
rect 554958 5216 554964 5228
rect 406896 5188 554964 5216
rect 406896 5176 406902 5188
rect 554958 5176 554964 5188
rect 555016 5176 555022 5228
rect 132954 5108 132960 5160
rect 133012 5148 133018 5160
rect 274634 5148 274640 5160
rect 133012 5120 274640 5148
rect 133012 5108 133018 5120
rect 274634 5108 274640 5120
rect 274692 5108 274698 5160
rect 278314 5108 278320 5160
rect 278372 5148 278378 5160
rect 320358 5148 320364 5160
rect 278372 5120 320364 5148
rect 278372 5108 278378 5120
rect 320358 5108 320364 5120
rect 320416 5108 320422 5160
rect 359918 5108 359924 5160
rect 359976 5148 359982 5160
rect 403618 5148 403624 5160
rect 359976 5120 403624 5148
rect 359976 5108 359982 5120
rect 403618 5108 403624 5120
rect 403676 5108 403682 5160
rect 408310 5108 408316 5160
rect 408368 5148 408374 5160
rect 558546 5148 558552 5160
rect 408368 5120 558552 5148
rect 408368 5108 408374 5120
rect 558546 5108 558552 5120
rect 558604 5108 558610 5160
rect 129366 5040 129372 5092
rect 129424 5080 129430 5092
rect 274726 5080 274732 5092
rect 129424 5052 274732 5080
rect 129424 5040 129430 5052
rect 274726 5040 274732 5052
rect 274784 5040 274790 5092
rect 274818 5040 274824 5092
rect 274876 5080 274882 5092
rect 318886 5080 318892 5092
rect 274876 5052 318892 5080
rect 274876 5040 274882 5052
rect 318886 5040 318892 5052
rect 318944 5040 318950 5092
rect 361206 5040 361212 5092
rect 361264 5080 361270 5092
rect 406010 5080 406016 5092
rect 361264 5052 406016 5080
rect 361264 5040 361270 5052
rect 406010 5040 406016 5052
rect 406068 5040 406074 5092
rect 409598 5040 409604 5092
rect 409656 5040 409662 5092
rect 409690 5040 409696 5092
rect 409748 5080 409754 5092
rect 562042 5080 562048 5092
rect 409748 5052 562048 5080
rect 409748 5040 409754 5052
rect 562042 5040 562048 5052
rect 562100 5040 562106 5092
rect 7650 4972 7656 5024
rect 7708 5012 7714 5024
rect 236086 5012 236092 5024
rect 7708 4984 236092 5012
rect 7708 4972 7714 4984
rect 236086 4972 236092 4984
rect 236144 4972 236150 5024
rect 246390 4972 246396 5024
rect 246448 5012 246454 5024
rect 310514 5012 310520 5024
rect 246448 4984 310520 5012
rect 246448 4972 246454 4984
rect 310514 4972 310520 4984
rect 310572 4972 310578 5024
rect 361298 4972 361304 5024
rect 361356 5012 361362 5024
rect 407206 5012 407212 5024
rect 361356 4984 407212 5012
rect 361356 4972 361362 4984
rect 407206 4972 407212 4984
rect 407264 4972 407270 5024
rect 409616 5012 409644 5040
rect 565630 5012 565636 5024
rect 409616 4984 565636 5012
rect 565630 4972 565636 4984
rect 565688 4972 565694 5024
rect 2866 4904 2872 4956
rect 2924 4944 2930 4956
rect 234798 4944 234804 4956
rect 2924 4916 234804 4944
rect 2924 4904 2930 4916
rect 234798 4904 234804 4916
rect 234856 4904 234862 4956
rect 242894 4904 242900 4956
rect 242952 4944 242958 4956
rect 309134 4944 309140 4956
rect 242952 4916 309140 4944
rect 242952 4904 242958 4916
rect 309134 4904 309140 4916
rect 309192 4904 309198 4956
rect 361390 4904 361396 4956
rect 361448 4944 361454 4956
rect 409598 4944 409604 4956
rect 361448 4916 409604 4944
rect 361448 4904 361454 4916
rect 409598 4904 409604 4916
rect 409656 4904 409662 4956
rect 411070 4904 411076 4956
rect 411128 4944 411134 4956
rect 569126 4944 569132 4956
rect 411128 4916 569132 4944
rect 411128 4904 411134 4916
rect 569126 4904 569132 4916
rect 569184 4904 569190 4956
rect 1670 4836 1676 4888
rect 1728 4876 1734 4888
rect 234890 4876 234896 4888
rect 1728 4848 234896 4876
rect 1728 4836 1734 4848
rect 234890 4836 234896 4848
rect 234948 4836 234954 4888
rect 239306 4836 239312 4888
rect 239364 4876 239370 4888
rect 307754 4876 307760 4888
rect 239364 4848 307760 4876
rect 239364 4836 239370 4848
rect 307754 4836 307760 4848
rect 307812 4836 307818 4888
rect 362678 4836 362684 4888
rect 362736 4876 362742 4888
rect 410794 4876 410800 4888
rect 362736 4848 410800 4876
rect 362736 4836 362742 4848
rect 410794 4836 410800 4848
rect 410852 4836 410858 4888
rect 412358 4836 412364 4888
rect 412416 4876 412422 4888
rect 572714 4876 572720 4888
rect 412416 4848 572720 4876
rect 412416 4836 412422 4848
rect 572714 4836 572720 4848
rect 572772 4836 572778 4888
rect 566 4768 572 4820
rect 624 4808 630 4820
rect 234706 4808 234712 4820
rect 624 4780 234712 4808
rect 624 4768 630 4780
rect 234706 4768 234712 4780
rect 234764 4768 234770 4820
rect 235810 4768 235816 4820
rect 235868 4808 235874 4820
rect 306466 4808 306472 4820
rect 235868 4780 306472 4808
rect 235868 4768 235874 4780
rect 306466 4768 306472 4780
rect 306524 4768 306530 4820
rect 362770 4768 362776 4820
rect 362828 4808 362834 4820
rect 413094 4808 413100 4820
rect 362828 4780 413100 4808
rect 362828 4768 362834 4780
rect 413094 4768 413100 4780
rect 413152 4768 413158 4820
rect 413830 4768 413836 4820
rect 413888 4808 413894 4820
rect 576302 4808 576308 4820
rect 413888 4780 576308 4808
rect 413888 4768 413894 4780
rect 576302 4768 576308 4780
rect 576360 4768 576366 4820
rect 193214 4700 193220 4752
rect 193272 4740 193278 4752
rect 220078 4740 220084 4752
rect 193272 4712 220084 4740
rect 193272 4700 193278 4712
rect 220078 4700 220084 4712
rect 220136 4700 220142 4752
rect 221550 4700 221556 4752
rect 221608 4740 221614 4752
rect 302510 4740 302516 4752
rect 221608 4712 302516 4740
rect 221608 4700 221614 4712
rect 302510 4700 302516 4712
rect 302568 4700 302574 4752
rect 355870 4700 355876 4752
rect 355928 4740 355934 4752
rect 388254 4740 388260 4752
rect 355928 4712 388260 4740
rect 355928 4700 355934 4712
rect 388254 4700 388260 4712
rect 388312 4700 388318 4752
rect 401318 4700 401324 4752
rect 401376 4740 401382 4752
rect 537202 4740 537208 4752
rect 401376 4712 537208 4740
rect 401376 4700 401382 4712
rect 537202 4700 537208 4712
rect 537260 4700 537266 4752
rect 171962 4632 171968 4684
rect 172020 4672 172026 4684
rect 222838 4672 222844 4684
rect 172020 4644 222844 4672
rect 172020 4632 172026 4644
rect 222838 4632 222844 4644
rect 222896 4632 222902 4684
rect 225138 4632 225144 4684
rect 225196 4672 225202 4684
rect 303798 4672 303804 4684
rect 225196 4644 303804 4672
rect 225196 4632 225202 4644
rect 303798 4632 303804 4644
rect 303856 4632 303862 4684
rect 354490 4632 354496 4684
rect 354548 4672 354554 4684
rect 384758 4672 384764 4684
rect 354548 4644 384764 4672
rect 354548 4632 354554 4644
rect 384758 4632 384764 4644
rect 384816 4632 384822 4684
rect 399846 4632 399852 4684
rect 399904 4672 399910 4684
rect 533706 4672 533712 4684
rect 399904 4644 533712 4672
rect 399904 4632 399910 4644
rect 533706 4632 533712 4644
rect 533764 4632 533770 4684
rect 228726 4564 228732 4616
rect 228784 4604 228790 4616
rect 304994 4604 305000 4616
rect 228784 4576 305000 4604
rect 228784 4564 228790 4576
rect 304994 4564 305000 4576
rect 305052 4564 305058 4616
rect 353110 4564 353116 4616
rect 353168 4604 353174 4616
rect 381170 4604 381176 4616
rect 353168 4576 381176 4604
rect 353168 4564 353174 4576
rect 381170 4564 381176 4576
rect 381228 4564 381234 4616
rect 398650 4564 398656 4616
rect 398708 4604 398714 4616
rect 530118 4604 530124 4616
rect 398708 4576 530124 4604
rect 398708 4564 398714 4576
rect 530118 4564 530124 4576
rect 530176 4564 530182 4616
rect 232222 4496 232228 4548
rect 232280 4536 232286 4548
rect 306374 4536 306380 4548
rect 232280 4508 306380 4536
rect 232280 4496 232286 4508
rect 306374 4496 306380 4508
rect 306432 4496 306438 4548
rect 351730 4496 351736 4548
rect 351788 4536 351794 4548
rect 377674 4536 377680 4548
rect 351788 4508 377680 4536
rect 351788 4496 351794 4508
rect 377674 4496 377680 4508
rect 377732 4496 377738 4548
rect 398558 4496 398564 4548
rect 398616 4536 398622 4548
rect 526622 4536 526628 4548
rect 398616 4508 526628 4536
rect 398616 4496 398622 4508
rect 526622 4496 526628 4508
rect 526680 4496 526686 4548
rect 281902 4428 281908 4480
rect 281960 4468 281966 4480
rect 321738 4468 321744 4480
rect 281960 4440 321744 4468
rect 281960 4428 281966 4440
rect 321738 4428 321744 4440
rect 321796 4428 321802 4480
rect 350258 4428 350264 4480
rect 350316 4468 350322 4480
rect 374086 4468 374092 4480
rect 350316 4440 374092 4468
rect 350316 4428 350322 4440
rect 374086 4428 374092 4440
rect 374144 4428 374150 4480
rect 397086 4428 397092 4480
rect 397144 4468 397150 4480
rect 523034 4468 523040 4480
rect 397144 4440 523040 4468
rect 397144 4428 397150 4440
rect 523034 4428 523040 4440
rect 523092 4428 523098 4480
rect 285398 4360 285404 4412
rect 285456 4400 285462 4412
rect 323026 4400 323032 4412
rect 285456 4372 323032 4400
rect 285456 4360 285462 4372
rect 323026 4360 323032 4372
rect 323084 4360 323090 4412
rect 395798 4360 395804 4412
rect 395856 4400 395862 4412
rect 519538 4400 519544 4412
rect 395856 4372 519544 4400
rect 395856 4360 395862 4372
rect 519538 4360 519544 4372
rect 519596 4360 519602 4412
rect 288986 4292 288992 4344
rect 289044 4332 289050 4344
rect 323118 4332 323124 4344
rect 289044 4304 323124 4332
rect 289044 4292 289050 4304
rect 323118 4292 323124 4304
rect 323176 4292 323182 4344
rect 394418 4292 394424 4344
rect 394476 4332 394482 4344
rect 515950 4332 515956 4344
rect 394476 4304 515956 4332
rect 394476 4292 394482 4304
rect 515950 4292 515956 4304
rect 516008 4292 516014 4344
rect 200298 4224 200304 4276
rect 200356 4264 200362 4276
rect 208946 4264 208952 4276
rect 200356 4236 208952 4264
rect 200356 4224 200362 4236
rect 208946 4224 208952 4236
rect 209004 4224 209010 4276
rect 292574 4224 292580 4276
rect 292632 4264 292638 4276
rect 324590 4264 324596 4276
rect 292632 4236 324596 4264
rect 292632 4224 292638 4236
rect 324590 4224 324596 4236
rect 324648 4224 324654 4276
rect 332594 4224 332600 4276
rect 332652 4264 332658 4276
rect 332778 4264 332784 4276
rect 332652 4236 332784 4264
rect 332652 4224 332658 4236
rect 332778 4224 332784 4236
rect 332836 4224 332842 4276
rect 392946 4224 392952 4276
rect 393004 4264 393010 4276
rect 512454 4264 512460 4276
rect 393004 4236 512460 4264
rect 393004 4224 393010 4236
rect 512454 4224 512460 4236
rect 512512 4224 512518 4276
rect 143534 4156 143540 4208
rect 143592 4196 143598 4208
rect 144822 4196 144828 4208
rect 143592 4168 144828 4196
rect 143592 4156 143598 4168
rect 144822 4156 144828 4168
rect 144880 4156 144886 4208
rect 184934 4156 184940 4208
rect 184992 4196 184998 4208
rect 186130 4196 186136 4208
rect 184992 4168 186136 4196
rect 184992 4156 184998 4168
rect 186130 4156 186136 4168
rect 186188 4156 186194 4208
rect 201494 4156 201500 4208
rect 201552 4196 201558 4208
rect 202782 4196 202788 4208
rect 201552 4168 202788 4196
rect 201552 4156 201558 4168
rect 202782 4156 202788 4168
rect 202840 4156 202846 4208
rect 226334 4156 226340 4208
rect 226392 4196 226398 4208
rect 227622 4196 227628 4208
rect 226392 4168 227628 4196
rect 226392 4156 226398 4168
rect 227622 4156 227628 4168
rect 227680 4156 227686 4208
rect 388438 4156 388444 4208
rect 388496 4196 388502 4208
rect 393038 4196 393044 4208
rect 388496 4168 393044 4196
rect 388496 4156 388502 4168
rect 393038 4156 393044 4168
rect 393096 4156 393102 4208
rect 418798 4156 418804 4208
rect 418856 4196 418862 4208
rect 420178 4196 420184 4208
rect 418856 4168 420184 4196
rect 418856 4156 418862 4168
rect 420178 4156 420184 4168
rect 420236 4156 420242 4208
rect 11146 4088 11152 4140
rect 11204 4128 11210 4140
rect 18598 4128 18604 4140
rect 11204 4100 18604 4128
rect 11204 4088 11210 4100
rect 18598 4088 18604 4100
rect 18656 4088 18662 4140
rect 34790 4088 34796 4140
rect 34848 4128 34854 4140
rect 36538 4128 36544 4140
rect 34848 4100 36544 4128
rect 34848 4088 34854 4100
rect 36538 4088 36544 4100
rect 36596 4088 36602 4140
rect 259730 4128 259736 4140
rect 84166 4100 259736 4128
rect 82078 4020 82084 4072
rect 82136 4060 82142 4072
rect 84166 4060 84194 4100
rect 259730 4088 259736 4100
rect 259788 4088 259794 4140
rect 306742 4088 306748 4140
rect 306800 4128 306806 4140
rect 328546 4128 328552 4140
rect 306800 4100 328552 4128
rect 306800 4088 306806 4100
rect 328546 4088 328552 4100
rect 328604 4088 328610 4140
rect 343542 4088 343548 4140
rect 343600 4128 343606 4140
rect 350442 4128 350448 4140
rect 343600 4100 350448 4128
rect 343600 4088 343606 4100
rect 350442 4088 350448 4100
rect 350500 4088 350506 4140
rect 351822 4088 351828 4140
rect 351880 4128 351886 4140
rect 375282 4128 375288 4140
rect 351880 4100 375288 4128
rect 351880 4088 351886 4100
rect 375282 4088 375288 4100
rect 375340 4088 375346 4140
rect 402790 4088 402796 4140
rect 402848 4128 402854 4140
rect 534997 4131 535055 4137
rect 534997 4128 535009 4131
rect 402848 4100 535009 4128
rect 402848 4088 402854 4100
rect 534997 4097 535009 4100
rect 535043 4097 535055 4131
rect 534997 4091 535055 4097
rect 82136 4032 84194 4060
rect 84381 4063 84439 4069
rect 82136 4020 82142 4032
rect 84381 4029 84393 4063
rect 84427 4060 84439 4063
rect 258166 4060 258172 4072
rect 84427 4032 258172 4060
rect 84427 4029 84439 4032
rect 84381 4023 84439 4029
rect 258166 4020 258172 4032
rect 258224 4020 258230 4072
rect 309042 4020 309048 4072
rect 309100 4060 309106 4072
rect 330110 4060 330116 4072
rect 309100 4032 330116 4060
rect 309100 4020 309106 4032
rect 330110 4020 330116 4032
rect 330168 4020 330174 4072
rect 332686 4020 332692 4072
rect 332744 4060 332750 4072
rect 335998 4060 336004 4072
rect 332744 4032 336004 4060
rect 332744 4020 332750 4032
rect 335998 4020 336004 4032
rect 336056 4020 336062 4072
rect 343450 4020 343456 4072
rect 343508 4060 343514 4072
rect 348050 4060 348056 4072
rect 343508 4032 348056 4060
rect 343508 4020 343514 4032
rect 348050 4020 348056 4032
rect 348108 4020 348114 4072
rect 350350 4020 350356 4072
rect 350408 4060 350414 4072
rect 372890 4060 372896 4072
rect 350408 4032 372896 4060
rect 350408 4020 350414 4032
rect 372890 4020 372896 4032
rect 372948 4020 372954 4072
rect 402606 4020 402612 4072
rect 402664 4060 402670 4072
rect 543182 4060 543188 4072
rect 402664 4032 543188 4060
rect 402664 4020 402670 4032
rect 543182 4020 543188 4032
rect 543240 4020 543246 4072
rect 43070 3952 43076 4004
rect 43128 3992 43134 4004
rect 51718 3992 51724 4004
rect 43128 3964 51724 3992
rect 43128 3952 43134 3964
rect 51718 3952 51724 3964
rect 51776 3952 51782 4004
rect 53650 3952 53656 4004
rect 53708 3992 53714 4004
rect 57238 3992 57244 4004
rect 53708 3964 57244 3992
rect 53708 3952 53714 3964
rect 57238 3952 57244 3964
rect 57296 3952 57302 4004
rect 74994 3952 75000 4004
rect 75052 3992 75058 4004
rect 258074 3992 258080 4004
rect 75052 3964 258080 3992
rect 75052 3952 75058 3964
rect 258074 3952 258080 3964
rect 258132 3952 258138 4004
rect 305546 3952 305552 4004
rect 305604 3992 305610 4004
rect 328730 3992 328736 4004
rect 305604 3964 328736 3992
rect 305604 3952 305610 3964
rect 328730 3952 328736 3964
rect 328788 3952 328794 4004
rect 329190 3952 329196 4004
rect 329248 3992 329254 4004
rect 335538 3992 335544 4004
rect 329248 3964 335544 3992
rect 329248 3952 329254 3964
rect 335538 3952 335544 3964
rect 335596 3952 335602 4004
rect 342162 3952 342168 4004
rect 342220 3992 342226 4004
rect 346946 3992 346952 4004
rect 342220 3964 346952 3992
rect 342220 3952 342226 3964
rect 346946 3952 346952 3964
rect 347004 3952 347010 4004
rect 353202 3952 353208 4004
rect 353260 3992 353266 4004
rect 379974 3992 379980 4004
rect 353260 3964 379980 3992
rect 353260 3952 353266 3964
rect 379974 3952 379980 3964
rect 380032 3952 380038 4004
rect 404262 3952 404268 4004
rect 404320 3992 404326 4004
rect 546678 3992 546684 4004
rect 404320 3964 546684 3992
rect 404320 3952 404326 3964
rect 546678 3952 546684 3964
rect 546736 3952 546742 4004
rect 38378 3884 38384 3936
rect 38436 3924 38442 3936
rect 47578 3924 47584 3936
rect 38436 3896 47584 3924
rect 38436 3884 38442 3896
rect 47578 3884 47584 3896
rect 47636 3884 47642 3936
rect 50154 3884 50160 3936
rect 50212 3924 50218 3936
rect 68278 3924 68284 3936
rect 50212 3896 68284 3924
rect 50212 3884 50218 3896
rect 68278 3884 68284 3896
rect 68336 3884 68342 3936
rect 71498 3884 71504 3936
rect 71556 3924 71562 3936
rect 256694 3924 256700 3936
rect 71556 3896 256700 3924
rect 71556 3884 71562 3896
rect 256694 3884 256700 3896
rect 256752 3884 256758 3936
rect 301958 3884 301964 3936
rect 302016 3924 302022 3936
rect 318061 3927 318119 3933
rect 318061 3924 318073 3927
rect 302016 3896 318073 3924
rect 302016 3884 302022 3896
rect 318061 3893 318073 3896
rect 318107 3893 318119 3927
rect 318061 3887 318119 3893
rect 318153 3927 318211 3933
rect 318153 3893 318165 3927
rect 318199 3924 318211 3927
rect 320361 3927 320419 3933
rect 320361 3924 320373 3927
rect 318199 3896 320373 3924
rect 318199 3893 318211 3896
rect 318153 3887 318211 3893
rect 320361 3893 320373 3896
rect 320407 3893 320419 3927
rect 325786 3924 325792 3936
rect 320361 3887 320419 3893
rect 320836 3896 325792 3924
rect 5258 3816 5264 3868
rect 5316 3856 5322 3868
rect 7558 3856 7564 3868
rect 5316 3828 7564 3856
rect 5316 3816 5322 3828
rect 7558 3816 7564 3828
rect 7616 3816 7622 3868
rect 41874 3816 41880 3868
rect 41932 3856 41938 3868
rect 54478 3856 54484 3868
rect 41932 3828 54484 3856
rect 41932 3816 41938 3828
rect 54478 3816 54484 3828
rect 54536 3816 54542 3868
rect 67910 3816 67916 3868
rect 67968 3856 67974 3868
rect 255314 3856 255320 3868
rect 67968 3828 255320 3856
rect 67968 3816 67974 3828
rect 255314 3816 255320 3828
rect 255372 3816 255378 3868
rect 297266 3816 297272 3868
rect 297324 3856 297330 3868
rect 320836 3856 320864 3896
rect 325786 3884 325792 3896
rect 325844 3884 325850 3936
rect 326798 3884 326804 3936
rect 326856 3924 326862 3936
rect 335630 3924 335636 3936
rect 326856 3896 335636 3924
rect 326856 3884 326862 3896
rect 335630 3884 335636 3896
rect 335688 3884 335694 3936
rect 344278 3884 344284 3936
rect 344336 3924 344342 3936
rect 351638 3924 351644 3936
rect 344336 3896 351644 3924
rect 344336 3884 344342 3896
rect 351638 3884 351644 3896
rect 351696 3884 351702 3936
rect 354582 3884 354588 3936
rect 354640 3924 354646 3936
rect 387150 3924 387156 3936
rect 354640 3896 387156 3924
rect 354640 3884 354646 3896
rect 387150 3884 387156 3896
rect 387208 3884 387214 3936
rect 405642 3884 405648 3936
rect 405700 3924 405706 3936
rect 550266 3924 550272 3936
rect 405700 3896 550272 3924
rect 405700 3884 405706 3896
rect 550266 3884 550272 3896
rect 550324 3884 550330 3936
rect 297324 3828 320864 3856
rect 297324 3816 297330 3828
rect 320910 3816 320916 3868
rect 320968 3856 320974 3868
rect 329098 3856 329104 3868
rect 320968 3828 329104 3856
rect 320968 3816 320974 3828
rect 329098 3816 329104 3828
rect 329156 3816 329162 3868
rect 333882 3816 333888 3868
rect 333940 3856 333946 3868
rect 336918 3856 336924 3868
rect 333940 3828 336924 3856
rect 333940 3816 333946 3828
rect 336918 3816 336924 3828
rect 336976 3816 336982 3868
rect 345750 3816 345756 3868
rect 345808 3856 345814 3868
rect 356330 3856 356336 3868
rect 345808 3828 356336 3856
rect 345808 3816 345814 3828
rect 356330 3816 356336 3828
rect 356388 3816 356394 3868
rect 357342 3816 357348 3868
rect 357400 3856 357406 3868
rect 358909 3859 358967 3865
rect 357400 3828 358860 3856
rect 357400 3816 357406 3828
rect 35986 3748 35992 3800
rect 36044 3788 36050 3800
rect 50338 3788 50344 3800
rect 36044 3760 50344 3788
rect 36044 3748 36050 3760
rect 50338 3748 50344 3760
rect 50396 3748 50402 3800
rect 64322 3748 64328 3800
rect 64380 3788 64386 3800
rect 253934 3788 253940 3800
rect 64380 3760 253940 3788
rect 64380 3748 64386 3760
rect 253934 3748 253940 3760
rect 253992 3748 253998 3800
rect 293678 3748 293684 3800
rect 293736 3788 293742 3800
rect 317969 3791 318027 3797
rect 317969 3788 317981 3791
rect 293736 3760 317981 3788
rect 293736 3748 293742 3760
rect 317969 3757 317981 3760
rect 318015 3757 318027 3791
rect 317969 3751 318027 3757
rect 318061 3791 318119 3797
rect 318061 3757 318073 3791
rect 318107 3788 318119 3791
rect 327258 3788 327264 3800
rect 318107 3760 327264 3788
rect 318107 3757 318119 3760
rect 318061 3751 318119 3757
rect 327258 3748 327264 3760
rect 327316 3748 327322 3800
rect 329009 3791 329067 3797
rect 329009 3757 329021 3791
rect 329055 3788 329067 3791
rect 334066 3788 334072 3800
rect 329055 3760 334072 3788
rect 329055 3757 329067 3760
rect 329009 3751 329067 3757
rect 334066 3748 334072 3760
rect 334124 3748 334130 3800
rect 343358 3748 343364 3800
rect 343416 3788 343422 3800
rect 349246 3788 349252 3800
rect 343416 3760 349252 3788
rect 343416 3748 343422 3760
rect 349246 3748 349252 3760
rect 349304 3748 349310 3800
rect 355962 3748 355968 3800
rect 356020 3788 356026 3800
rect 358633 3791 358691 3797
rect 358633 3788 358645 3791
rect 356020 3760 358645 3788
rect 356020 3748 356026 3760
rect 358633 3757 358645 3760
rect 358679 3757 358691 3791
rect 358633 3751 358691 3757
rect 358722 3748 358728 3800
rect 358780 3748 358786 3800
rect 358832 3788 358860 3828
rect 358909 3825 358921 3859
rect 358955 3856 358967 3859
rect 390646 3856 390652 3868
rect 358955 3828 390652 3856
rect 358955 3825 358967 3828
rect 358909 3819 358967 3825
rect 390646 3816 390652 3828
rect 390704 3816 390710 3868
rect 406930 3816 406936 3868
rect 406988 3856 406994 3868
rect 553762 3856 553768 3868
rect 406988 3828 553768 3856
rect 406988 3816 406994 3828
rect 553762 3816 553768 3828
rect 553820 3816 553826 3868
rect 394234 3788 394240 3800
rect 358832 3760 394240 3788
rect 394234 3748 394240 3760
rect 394292 3748 394298 3800
rect 407022 3748 407028 3800
rect 407080 3788 407086 3800
rect 557350 3788 557356 3800
rect 407080 3760 557356 3788
rect 407080 3748 407086 3760
rect 557350 3748 557356 3760
rect 557408 3748 557414 3800
rect 23014 3680 23020 3732
rect 23072 3720 23078 3732
rect 39298 3720 39304 3732
rect 23072 3692 39304 3720
rect 23072 3680 23078 3692
rect 39298 3680 39304 3692
rect 39356 3680 39362 3732
rect 43438 3720 43444 3732
rect 39500 3692 43444 3720
rect 20622 3612 20628 3664
rect 20680 3652 20686 3664
rect 39500 3652 39528 3692
rect 43438 3680 43444 3692
rect 43496 3680 43502 3732
rect 45370 3680 45376 3732
rect 45428 3720 45434 3732
rect 58618 3720 58624 3732
rect 45428 3692 58624 3720
rect 45428 3680 45434 3692
rect 58618 3680 58624 3692
rect 58676 3680 58682 3732
rect 60826 3680 60832 3732
rect 60884 3720 60890 3732
rect 252830 3720 252836 3732
rect 60884 3692 252836 3720
rect 60884 3680 60890 3692
rect 252830 3680 252836 3692
rect 252888 3680 252894 3732
rect 291378 3680 291384 3732
rect 291436 3720 291442 3732
rect 324314 3720 324320 3732
rect 291436 3692 324320 3720
rect 291436 3680 291442 3692
rect 324314 3680 324320 3692
rect 324372 3680 324378 3732
rect 324406 3680 324412 3732
rect 324464 3720 324470 3732
rect 334158 3720 334164 3732
rect 324464 3692 334164 3720
rect 324464 3680 324470 3692
rect 334158 3680 334164 3692
rect 334216 3680 334222 3732
rect 346302 3680 346308 3732
rect 346360 3720 346366 3732
rect 358740 3720 358768 3748
rect 397730 3720 397736 3732
rect 346360 3692 353156 3720
rect 358740 3692 397736 3720
rect 346360 3680 346366 3692
rect 20680 3624 39528 3652
rect 20680 3612 20686 3624
rect 39574 3612 39580 3664
rect 39632 3652 39638 3664
rect 53929 3655 53987 3661
rect 39632 3624 53880 3652
rect 39632 3612 39638 3624
rect 18230 3544 18236 3596
rect 18288 3584 18294 3596
rect 18288 3556 26234 3584
rect 18288 3544 18294 3556
rect 26206 3516 26234 3556
rect 28902 3544 28908 3596
rect 28960 3584 28966 3596
rect 35158 3584 35164 3596
rect 28960 3556 35164 3584
rect 28960 3544 28966 3556
rect 35158 3544 35164 3556
rect 35216 3544 35222 3596
rect 40678 3544 40684 3596
rect 40736 3584 40742 3596
rect 41322 3584 41328 3596
rect 40736 3556 41328 3584
rect 40736 3544 40742 3556
rect 41322 3544 41328 3556
rect 41380 3544 41386 3596
rect 48958 3544 48964 3596
rect 49016 3584 49022 3596
rect 49602 3584 49608 3596
rect 49016 3556 49608 3584
rect 49016 3544 49022 3556
rect 49602 3544 49608 3556
rect 49660 3544 49666 3596
rect 52546 3544 52552 3596
rect 52604 3584 52610 3596
rect 53742 3584 53748 3596
rect 52604 3556 53748 3584
rect 52604 3544 52610 3556
rect 53742 3544 53748 3556
rect 53800 3544 53806 3596
rect 53852 3584 53880 3624
rect 53929 3621 53941 3655
rect 53975 3652 53987 3655
rect 248690 3652 248696 3664
rect 53975 3624 248696 3652
rect 53975 3621 53987 3624
rect 53929 3615 53987 3621
rect 248690 3612 248696 3624
rect 248748 3612 248754 3664
rect 284294 3612 284300 3664
rect 284352 3652 284358 3664
rect 321830 3652 321836 3664
rect 284352 3624 321836 3652
rect 284352 3612 284358 3624
rect 321830 3612 321836 3624
rect 321888 3612 321894 3664
rect 324498 3652 324504 3664
rect 321940 3624 324504 3652
rect 247218 3584 247224 3596
rect 53852 3556 247224 3584
rect 247218 3544 247224 3556
rect 247276 3544 247282 3596
rect 279510 3544 279516 3596
rect 279568 3584 279574 3596
rect 279568 3556 281580 3584
rect 279568 3544 279574 3556
rect 32306 3516 32312 3528
rect 26206 3488 32312 3516
rect 32306 3476 32312 3488
rect 32364 3476 32370 3528
rect 32398 3476 32404 3528
rect 32456 3516 32462 3528
rect 244458 3516 244464 3528
rect 32456 3488 244464 3516
rect 32456 3476 32462 3488
rect 244458 3476 244464 3488
rect 244516 3476 244522 3528
rect 249978 3476 249984 3528
rect 250036 3516 250042 3528
rect 251082 3516 251088 3528
rect 250036 3488 251088 3516
rect 250036 3476 250042 3488
rect 251082 3476 251088 3488
rect 251140 3476 251146 3528
rect 255866 3476 255872 3528
rect 255924 3516 255930 3528
rect 256602 3516 256608 3528
rect 255924 3488 256608 3516
rect 255924 3476 255930 3488
rect 256602 3476 256608 3488
rect 256660 3476 256666 3528
rect 262950 3476 262956 3528
rect 263008 3516 263014 3528
rect 263502 3516 263508 3528
rect 263008 3488 263508 3516
rect 263008 3476 263014 3488
rect 263502 3476 263508 3488
rect 263560 3476 263566 3528
rect 264146 3476 264152 3528
rect 264204 3516 264210 3528
rect 264882 3516 264888 3528
rect 264204 3488 264888 3516
rect 264204 3476 264210 3488
rect 264882 3476 264888 3488
rect 264940 3476 264946 3528
rect 266538 3476 266544 3528
rect 266596 3516 266602 3528
rect 267642 3516 267648 3528
rect 266596 3488 267648 3516
rect 266596 3476 266602 3488
rect 267642 3476 267648 3488
rect 267700 3476 267706 3528
rect 271230 3476 271236 3528
rect 271288 3516 271294 3528
rect 271782 3516 271788 3528
rect 271288 3488 271788 3516
rect 271288 3476 271294 3488
rect 271782 3476 271788 3488
rect 271840 3476 271846 3528
rect 273622 3476 273628 3528
rect 273680 3516 273686 3528
rect 274542 3516 274548 3528
rect 273680 3488 274548 3516
rect 273680 3476 273686 3488
rect 274542 3476 274548 3488
rect 274600 3476 274606 3528
rect 276014 3476 276020 3528
rect 276072 3516 276078 3528
rect 277302 3516 277308 3528
rect 276072 3488 277308 3516
rect 276072 3476 276078 3488
rect 277302 3476 277308 3488
rect 277360 3476 277366 3528
rect 280706 3476 280712 3528
rect 280764 3516 280770 3528
rect 281442 3516 281448 3528
rect 280764 3488 281448 3516
rect 280764 3476 280770 3488
rect 281442 3476 281448 3488
rect 281500 3476 281506 3528
rect 281552 3516 281580 3556
rect 286594 3544 286600 3596
rect 286652 3584 286658 3596
rect 317877 3587 317935 3593
rect 317877 3584 317889 3587
rect 286652 3556 317889 3584
rect 286652 3544 286658 3556
rect 317877 3553 317889 3556
rect 317923 3553 317935 3587
rect 317877 3547 317935 3553
rect 317969 3587 318027 3593
rect 317969 3553 317981 3587
rect 318015 3584 318027 3587
rect 321940 3584 321968 3624
rect 324498 3612 324504 3624
rect 324556 3612 324562 3664
rect 325602 3612 325608 3664
rect 325660 3652 325666 3664
rect 335446 3652 335452 3664
rect 325660 3624 335452 3652
rect 325660 3612 325666 3624
rect 335446 3612 335452 3624
rect 335504 3612 335510 3664
rect 347130 3612 347136 3664
rect 347188 3652 347194 3664
rect 353128 3652 353156 3692
rect 397730 3680 397736 3692
rect 397788 3680 397794 3732
rect 408402 3680 408408 3732
rect 408460 3720 408466 3732
rect 560846 3720 560852 3732
rect 408460 3692 560852 3720
rect 408460 3680 408466 3692
rect 560846 3680 560852 3692
rect 560904 3680 560910 3732
rect 358722 3652 358728 3664
rect 347188 3624 353064 3652
rect 353128 3624 358728 3652
rect 347188 3612 347194 3624
rect 323210 3584 323216 3596
rect 318015 3556 321968 3584
rect 322032 3556 323216 3584
rect 318015 3553 318027 3556
rect 317969 3547 318027 3553
rect 320266 3516 320272 3528
rect 281552 3488 320272 3516
rect 320266 3476 320272 3488
rect 320324 3476 320330 3528
rect 320361 3519 320419 3525
rect 320361 3485 320373 3519
rect 320407 3516 320419 3519
rect 322032 3516 322060 3556
rect 323210 3544 323216 3556
rect 323268 3544 323274 3596
rect 323302 3544 323308 3596
rect 323360 3584 323366 3596
rect 329009 3587 329067 3593
rect 329009 3584 329021 3587
rect 323360 3556 329021 3584
rect 323360 3544 323366 3556
rect 329009 3553 329021 3556
rect 329055 3553 329067 3587
rect 329009 3547 329067 3553
rect 329193 3587 329251 3593
rect 329193 3553 329205 3587
rect 329239 3584 329251 3587
rect 332594 3584 332600 3596
rect 329239 3556 332600 3584
rect 329239 3553 329251 3556
rect 329193 3547 329251 3553
rect 332594 3544 332600 3556
rect 332652 3544 332658 3596
rect 342070 3544 342076 3596
rect 342128 3584 342134 3596
rect 344554 3584 344560 3596
rect 342128 3556 344560 3584
rect 342128 3544 342134 3556
rect 344554 3544 344560 3556
rect 344612 3544 344618 3596
rect 347590 3544 347596 3596
rect 347648 3584 347654 3596
rect 353036 3584 353064 3624
rect 358722 3612 358728 3624
rect 358780 3612 358786 3664
rect 360010 3612 360016 3664
rect 360068 3652 360074 3664
rect 401318 3652 401324 3664
rect 360068 3624 401324 3652
rect 360068 3612 360074 3624
rect 401318 3612 401324 3624
rect 401376 3612 401382 3664
rect 409782 3612 409788 3664
rect 409840 3652 409846 3664
rect 564434 3652 564440 3664
rect 409840 3624 564440 3652
rect 409840 3612 409846 3624
rect 564434 3612 564440 3624
rect 564492 3612 564498 3664
rect 359918 3584 359924 3596
rect 347648 3556 352972 3584
rect 353036 3556 359924 3584
rect 347648 3544 347654 3556
rect 320407 3488 322060 3516
rect 320407 3485 320419 3488
rect 320361 3479 320419 3485
rect 322106 3476 322112 3528
rect 322164 3516 322170 3528
rect 322164 3488 330064 3516
rect 322164 3476 322170 3488
rect 13538 3408 13544 3460
rect 13596 3448 13602 3460
rect 22738 3448 22744 3460
rect 13596 3420 22744 3448
rect 13596 3408 13602 3420
rect 22738 3408 22744 3420
rect 22796 3408 22802 3460
rect 25314 3408 25320 3460
rect 25372 3448 25378 3460
rect 241606 3448 241612 3460
rect 25372 3420 241612 3448
rect 25372 3408 25378 3420
rect 241606 3408 241612 3420
rect 241664 3408 241670 3460
rect 267734 3408 267740 3460
rect 267792 3448 267798 3460
rect 269022 3448 269028 3460
rect 267792 3420 269028 3448
rect 267792 3408 267798 3420
rect 269022 3408 269028 3420
rect 269080 3408 269086 3460
rect 272426 3408 272432 3460
rect 272484 3448 272490 3460
rect 318978 3448 318984 3460
rect 272484 3420 318984 3448
rect 272484 3408 272490 3420
rect 318978 3408 318984 3420
rect 319036 3408 319042 3460
rect 319714 3408 319720 3460
rect 319772 3448 319778 3460
rect 329193 3451 329251 3457
rect 329193 3448 329205 3451
rect 319772 3420 329205 3448
rect 319772 3408 319778 3420
rect 329193 3417 329205 3420
rect 329239 3417 329251 3451
rect 329193 3411 329251 3417
rect 19426 3340 19432 3392
rect 19484 3380 19490 3392
rect 25498 3380 25504 3392
rect 19484 3352 25504 3380
rect 19484 3340 19490 3352
rect 25498 3340 25504 3352
rect 25556 3340 25562 3392
rect 31294 3340 31300 3392
rect 31352 3380 31358 3392
rect 33778 3380 33784 3392
rect 31352 3352 33784 3380
rect 31352 3340 31358 3352
rect 33778 3340 33784 3352
rect 33836 3340 33842 3392
rect 44266 3340 44272 3392
rect 44324 3380 44330 3392
rect 45462 3380 45468 3392
rect 44324 3352 45468 3380
rect 44324 3340 44330 3352
rect 45462 3340 45468 3352
rect 45520 3340 45526 3392
rect 46658 3340 46664 3392
rect 46716 3380 46722 3392
rect 53929 3383 53987 3389
rect 53929 3380 53941 3383
rect 46716 3352 53941 3380
rect 46716 3340 46722 3352
rect 53929 3349 53941 3352
rect 53975 3349 53987 3383
rect 53929 3343 53987 3349
rect 56042 3340 56048 3392
rect 56100 3380 56106 3392
rect 56502 3380 56508 3392
rect 56100 3352 56508 3380
rect 56100 3340 56106 3352
rect 56502 3340 56508 3352
rect 56560 3340 56566 3392
rect 59630 3340 59636 3392
rect 59688 3380 59694 3392
rect 60642 3380 60648 3392
rect 59688 3352 60648 3380
rect 59688 3340 59694 3352
rect 60642 3340 60648 3352
rect 60700 3340 60706 3392
rect 66714 3340 66720 3392
rect 66772 3380 66778 3392
rect 67542 3380 67548 3392
rect 66772 3352 67548 3380
rect 66772 3340 66778 3352
rect 67542 3340 67548 3352
rect 67600 3340 67606 3392
rect 73798 3340 73804 3392
rect 73856 3380 73862 3392
rect 74442 3380 74448 3392
rect 73856 3352 74448 3380
rect 73856 3340 73862 3352
rect 74442 3340 74448 3352
rect 74500 3340 74506 3392
rect 77386 3340 77392 3392
rect 77444 3380 77450 3392
rect 78582 3380 78588 3392
rect 77444 3352 78588 3380
rect 77444 3340 77450 3352
rect 78582 3340 78588 3352
rect 78640 3340 78646 3392
rect 80882 3340 80888 3392
rect 80940 3380 80946 3392
rect 81342 3380 81348 3392
rect 80940 3352 81348 3380
rect 80940 3340 80946 3352
rect 81342 3340 81348 3352
rect 81400 3340 81406 3392
rect 84381 3383 84439 3389
rect 84381 3380 84393 3383
rect 81452 3352 84393 3380
rect 78582 3204 78588 3256
rect 78640 3244 78646 3256
rect 81452 3244 81480 3352
rect 84381 3349 84393 3352
rect 84427 3349 84439 3383
rect 84381 3343 84439 3349
rect 84470 3340 84476 3392
rect 84528 3380 84534 3392
rect 87598 3380 87604 3392
rect 84528 3352 87604 3380
rect 84528 3340 84534 3352
rect 87598 3340 87604 3352
rect 87656 3340 87662 3392
rect 90358 3340 90364 3392
rect 90416 3380 90422 3392
rect 91002 3380 91008 3392
rect 90416 3352 91008 3380
rect 90416 3340 90422 3352
rect 91002 3340 91008 3352
rect 91060 3340 91066 3392
rect 91554 3340 91560 3392
rect 91612 3380 91618 3392
rect 93118 3380 93124 3392
rect 91612 3352 93124 3380
rect 91612 3340 91618 3352
rect 93118 3340 93124 3352
rect 93176 3340 93182 3392
rect 261018 3380 261024 3392
rect 93826 3352 261024 3380
rect 83274 3272 83280 3324
rect 83332 3312 83338 3324
rect 84102 3312 84108 3324
rect 83332 3284 84108 3312
rect 83332 3272 83338 3284
rect 84102 3272 84108 3284
rect 84160 3272 84166 3324
rect 87966 3272 87972 3324
rect 88024 3312 88030 3324
rect 88978 3312 88984 3324
rect 88024 3284 88984 3312
rect 88024 3272 88030 3284
rect 88978 3272 88984 3284
rect 89036 3272 89042 3324
rect 93826 3312 93854 3352
rect 261018 3340 261024 3352
rect 261076 3340 261082 3392
rect 287790 3340 287796 3392
rect 287848 3380 287854 3392
rect 288342 3380 288348 3392
rect 287848 3352 288348 3380
rect 287848 3340 287854 3352
rect 288342 3340 288348 3352
rect 288400 3340 288406 3392
rect 296070 3340 296076 3392
rect 296128 3380 296134 3392
rect 296622 3380 296628 3392
rect 296128 3352 296628 3380
rect 296128 3340 296134 3352
rect 296622 3340 296628 3352
rect 296680 3340 296686 3392
rect 298462 3340 298468 3392
rect 298520 3380 298526 3392
rect 299382 3380 299388 3392
rect 298520 3352 299388 3380
rect 298520 3340 298526 3352
rect 299382 3340 299388 3352
rect 299440 3340 299446 3392
rect 307938 3340 307944 3392
rect 307996 3380 308002 3392
rect 329834 3380 329840 3392
rect 307996 3352 329840 3380
rect 307996 3340 308002 3352
rect 329834 3340 329840 3352
rect 329892 3340 329898 3392
rect 330036 3380 330064 3488
rect 331582 3476 331588 3528
rect 331640 3516 331646 3528
rect 332502 3516 332508 3528
rect 331640 3488 332508 3516
rect 331640 3476 331646 3488
rect 332502 3476 332508 3488
rect 332560 3476 332566 3528
rect 337470 3476 337476 3528
rect 337528 3516 337534 3528
rect 338114 3516 338120 3528
rect 337528 3488 338120 3516
rect 337528 3476 337534 3488
rect 338114 3476 338120 3488
rect 338172 3476 338178 3528
rect 345658 3476 345664 3528
rect 345716 3516 345722 3528
rect 352834 3516 352840 3528
rect 345716 3488 352840 3516
rect 345716 3476 345722 3488
rect 352834 3476 352840 3488
rect 352892 3476 352898 3528
rect 352944 3516 352972 3556
rect 359918 3544 359924 3556
rect 359976 3544 359982 3596
rect 360102 3544 360108 3596
rect 360160 3584 360166 3596
rect 404814 3584 404820 3596
rect 360160 3556 404820 3584
rect 360160 3544 360166 3556
rect 404814 3544 404820 3556
rect 404872 3544 404878 3596
rect 411162 3544 411168 3596
rect 411220 3584 411226 3596
rect 568022 3584 568028 3596
rect 411220 3556 568028 3584
rect 411220 3544 411226 3556
rect 568022 3544 568028 3556
rect 568080 3544 568086 3596
rect 361114 3516 361120 3528
rect 352944 3488 361120 3516
rect 361114 3476 361120 3488
rect 361172 3476 361178 3528
rect 361482 3476 361488 3528
rect 361540 3516 361546 3528
rect 408402 3516 408408 3528
rect 361540 3488 408408 3516
rect 361540 3476 361546 3488
rect 408402 3476 408408 3488
rect 408460 3476 408466 3528
rect 412542 3476 412548 3528
rect 412600 3516 412606 3528
rect 571518 3516 571524 3528
rect 412600 3488 571524 3516
rect 412600 3476 412606 3488
rect 571518 3476 571524 3488
rect 571576 3476 571582 3528
rect 330386 3408 330392 3460
rect 330444 3448 330450 3460
rect 333238 3448 333244 3460
rect 330444 3420 333244 3448
rect 330444 3408 330450 3420
rect 333238 3408 333244 3420
rect 333296 3408 333302 3460
rect 335078 3408 335084 3460
rect 335136 3448 335142 3460
rect 338206 3448 338212 3460
rect 335136 3420 338212 3448
rect 335136 3408 335142 3420
rect 338206 3408 338212 3420
rect 338264 3408 338270 3460
rect 347682 3408 347688 3460
rect 347740 3448 347746 3460
rect 362310 3448 362316 3460
rect 347740 3420 362316 3448
rect 347740 3408 347746 3420
rect 362310 3408 362316 3420
rect 362368 3408 362374 3460
rect 362862 3408 362868 3460
rect 362920 3448 362926 3460
rect 411898 3448 411904 3460
rect 362920 3420 411904 3448
rect 362920 3408 362926 3420
rect 411898 3408 411904 3420
rect 411956 3408 411962 3460
rect 412450 3408 412456 3460
rect 412508 3448 412514 3460
rect 575106 3448 575112 3460
rect 412508 3420 575112 3448
rect 412508 3408 412514 3420
rect 575106 3408 575112 3420
rect 575164 3408 575170 3460
rect 334342 3380 334348 3392
rect 330036 3352 334348 3380
rect 334342 3340 334348 3352
rect 334400 3340 334406 3392
rect 350534 3340 350540 3392
rect 350592 3380 350598 3392
rect 371694 3380 371700 3392
rect 350592 3352 371700 3380
rect 350592 3340 350598 3352
rect 371694 3340 371700 3352
rect 371752 3340 371758 3392
rect 382182 3340 382188 3392
rect 382240 3380 382246 3392
rect 475746 3380 475752 3392
rect 382240 3352 475752 3380
rect 382240 3340 382246 3352
rect 475746 3340 475752 3352
rect 475804 3340 475810 3392
rect 481634 3340 481640 3392
rect 481692 3380 481698 3392
rect 482830 3380 482836 3392
rect 481692 3352 482836 3380
rect 481692 3340 481698 3352
rect 482830 3340 482836 3352
rect 482888 3340 482894 3392
rect 489178 3340 489184 3392
rect 489236 3380 489242 3392
rect 489914 3380 489920 3392
rect 489236 3352 489920 3380
rect 489236 3340 489242 3352
rect 489914 3340 489920 3352
rect 489972 3340 489978 3392
rect 499546 3352 528554 3380
rect 89732 3284 93854 3312
rect 78640 3216 81480 3244
rect 78640 3204 78646 3216
rect 85666 3204 85672 3256
rect 85724 3244 85730 3256
rect 89732 3244 89760 3284
rect 93946 3272 93952 3324
rect 94004 3312 94010 3324
rect 95050 3312 95056 3324
rect 94004 3284 95056 3312
rect 94004 3272 94010 3284
rect 95050 3272 95056 3284
rect 95108 3272 95114 3324
rect 97442 3272 97448 3324
rect 97500 3312 97506 3324
rect 97902 3312 97908 3324
rect 97500 3284 97908 3312
rect 97500 3272 97506 3284
rect 97902 3272 97908 3284
rect 97960 3272 97966 3324
rect 98638 3272 98644 3324
rect 98696 3312 98702 3324
rect 99282 3312 99288 3324
rect 98696 3284 99288 3312
rect 98696 3272 98702 3284
rect 99282 3272 99288 3284
rect 99340 3272 99346 3324
rect 101030 3272 101036 3324
rect 101088 3312 101094 3324
rect 102042 3312 102048 3324
rect 101088 3284 102048 3312
rect 101088 3272 101094 3284
rect 102042 3272 102048 3284
rect 102100 3272 102106 3324
rect 102137 3315 102195 3321
rect 102137 3281 102149 3315
rect 102183 3312 102195 3315
rect 262490 3312 262496 3324
rect 102183 3284 262496 3312
rect 102183 3281 102195 3284
rect 102137 3275 102195 3281
rect 262490 3272 262496 3284
rect 262548 3272 262554 3324
rect 310238 3272 310244 3324
rect 310296 3312 310302 3324
rect 330018 3312 330024 3324
rect 310296 3284 330024 3312
rect 310296 3272 310302 3284
rect 330018 3272 330024 3284
rect 330076 3272 330082 3324
rect 348970 3272 348976 3324
rect 349028 3312 349034 3324
rect 369394 3312 369400 3324
rect 349028 3284 369400 3312
rect 349028 3272 349034 3284
rect 369394 3272 369400 3284
rect 369452 3272 369458 3324
rect 380802 3272 380808 3324
rect 380860 3312 380866 3324
rect 468662 3312 468668 3324
rect 380860 3284 468668 3312
rect 380860 3272 380866 3284
rect 468662 3272 468668 3284
rect 468720 3272 468726 3324
rect 485038 3272 485044 3324
rect 485096 3312 485102 3324
rect 499546 3312 499574 3352
rect 485096 3284 499574 3312
rect 485096 3272 485102 3284
rect 502978 3272 502984 3324
rect 503036 3312 503042 3324
rect 504174 3312 504180 3324
rect 503036 3284 504180 3312
rect 503036 3272 503042 3284
rect 504174 3272 504180 3284
rect 504232 3272 504238 3324
rect 506474 3272 506480 3324
rect 506532 3312 506538 3324
rect 507670 3312 507676 3324
rect 506532 3284 507676 3312
rect 506532 3272 506538 3284
rect 507670 3272 507676 3284
rect 507728 3272 507734 3324
rect 515398 3272 515404 3324
rect 515456 3312 515462 3324
rect 517146 3312 517152 3324
rect 515456 3284 517152 3312
rect 515456 3272 515462 3284
rect 517146 3272 517152 3284
rect 517204 3272 517210 3324
rect 519630 3272 519636 3324
rect 519688 3312 519694 3324
rect 521838 3312 521844 3324
rect 519688 3284 521844 3312
rect 519688 3272 519694 3284
rect 521838 3272 521844 3284
rect 521896 3272 521902 3324
rect 522298 3272 522304 3324
rect 522356 3312 522362 3324
rect 524230 3312 524236 3324
rect 522356 3284 524236 3312
rect 522356 3272 522362 3284
rect 524230 3272 524236 3284
rect 524288 3272 524294 3324
rect 528526 3312 528554 3352
rect 530578 3340 530584 3392
rect 530636 3380 530642 3392
rect 531314 3380 531320 3392
rect 530636 3352 531320 3380
rect 530636 3340 530642 3352
rect 531314 3340 531320 3352
rect 531372 3340 531378 3392
rect 533338 3340 533344 3392
rect 533396 3380 533402 3392
rect 534902 3380 534908 3392
rect 533396 3352 534908 3380
rect 533396 3340 533402 3352
rect 534902 3340 534908 3352
rect 534960 3340 534966 3392
rect 534997 3383 535055 3389
rect 534997 3349 535009 3383
rect 535043 3380 535055 3383
rect 539594 3380 539600 3392
rect 535043 3352 539600 3380
rect 535043 3349 535055 3352
rect 534997 3343 535055 3349
rect 539594 3340 539600 3352
rect 539652 3340 539658 3392
rect 540238 3340 540244 3392
rect 540296 3380 540302 3392
rect 541986 3380 541992 3392
rect 540296 3352 541992 3380
rect 540296 3340 540302 3352
rect 541986 3340 541992 3352
rect 542044 3340 542050 3392
rect 532510 3312 532516 3324
rect 528526 3284 532516 3312
rect 532510 3272 532516 3284
rect 532568 3272 532574 3324
rect 85724 3216 89760 3244
rect 85724 3204 85730 3216
rect 92750 3204 92756 3256
rect 92808 3244 92814 3256
rect 262306 3244 262312 3256
rect 92808 3216 262312 3244
rect 92808 3204 92814 3216
rect 262306 3204 262312 3216
rect 262364 3204 262370 3256
rect 312630 3204 312636 3256
rect 312688 3244 312694 3256
rect 331398 3244 331404 3256
rect 312688 3216 331404 3244
rect 312688 3204 312694 3216
rect 331398 3204 331404 3216
rect 331456 3204 331462 3256
rect 349062 3204 349068 3256
rect 349120 3244 349126 3256
rect 365806 3244 365812 3256
rect 349120 3216 365812 3244
rect 349120 3204 349126 3216
rect 365806 3204 365812 3216
rect 365864 3204 365870 3256
rect 377766 3204 377772 3256
rect 377824 3244 377830 3256
rect 461578 3244 461584 3256
rect 377824 3216 461584 3244
rect 377824 3204 377830 3216
rect 461578 3204 461584 3216
rect 461636 3204 461642 3256
rect 526438 3204 526444 3256
rect 526496 3244 526502 3256
rect 527818 3244 527824 3256
rect 526496 3216 527824 3244
rect 526496 3204 526502 3216
rect 527818 3204 527824 3216
rect 527876 3204 527882 3256
rect 57238 3136 57244 3188
rect 57296 3176 57302 3188
rect 61378 3176 61384 3188
rect 57296 3148 61384 3176
rect 57296 3136 57302 3148
rect 61378 3136 61384 3148
rect 61436 3136 61442 3188
rect 89162 3136 89168 3188
rect 89220 3176 89226 3188
rect 102045 3179 102103 3185
rect 102045 3176 102057 3179
rect 89220 3148 102057 3176
rect 89220 3136 89226 3148
rect 102045 3145 102057 3148
rect 102091 3145 102103 3179
rect 263778 3176 263784 3188
rect 102045 3139 102103 3145
rect 102152 3148 263784 3176
rect 96246 3068 96252 3120
rect 96304 3108 96310 3120
rect 102152 3108 102180 3148
rect 263778 3136 263784 3148
rect 263836 3136 263842 3188
rect 311434 3136 311440 3188
rect 311492 3176 311498 3188
rect 329926 3176 329932 3188
rect 311492 3148 329932 3176
rect 311492 3136 311498 3148
rect 329926 3136 329932 3148
rect 329984 3136 329990 3188
rect 349798 3136 349804 3188
rect 349856 3176 349862 3188
rect 354217 3179 354275 3185
rect 349856 3148 354168 3176
rect 349856 3136 349862 3148
rect 96304 3080 102180 3108
rect 96304 3068 96310 3080
rect 102226 3068 102232 3120
rect 102284 3108 102290 3120
rect 104158 3108 104164 3120
rect 102284 3080 104164 3108
rect 102284 3068 102290 3080
rect 104158 3068 104164 3080
rect 104216 3068 104222 3120
rect 105722 3068 105728 3120
rect 105780 3108 105786 3120
rect 106182 3108 106188 3120
rect 105780 3080 106188 3108
rect 105780 3068 105786 3080
rect 106182 3068 106188 3080
rect 106240 3068 106246 3120
rect 106918 3068 106924 3120
rect 106976 3108 106982 3120
rect 107562 3108 107568 3120
rect 106976 3080 107568 3108
rect 106976 3068 106982 3080
rect 107562 3068 107568 3080
rect 107620 3068 107626 3120
rect 108114 3068 108120 3120
rect 108172 3108 108178 3120
rect 108942 3108 108948 3120
rect 108172 3080 108948 3108
rect 108172 3068 108178 3080
rect 108942 3068 108948 3080
rect 109000 3068 109006 3120
rect 109310 3068 109316 3120
rect 109368 3108 109374 3120
rect 111058 3108 111064 3120
rect 109368 3080 111064 3108
rect 109368 3068 109374 3080
rect 111058 3068 111064 3080
rect 111116 3068 111122 3120
rect 111153 3111 111211 3117
rect 111153 3077 111165 3111
rect 111199 3108 111211 3111
rect 265250 3108 265256 3120
rect 111199 3080 265256 3108
rect 111199 3077 111211 3080
rect 111153 3071 111211 3077
rect 265250 3068 265256 3080
rect 265308 3068 265314 3120
rect 313826 3068 313832 3120
rect 313884 3108 313890 3120
rect 331490 3108 331496 3120
rect 313884 3080 331496 3108
rect 313884 3068 313890 3080
rect 331490 3068 331496 3080
rect 331548 3068 331554 3120
rect 338666 3068 338672 3120
rect 338724 3108 338730 3120
rect 339586 3108 339592 3120
rect 338724 3080 339592 3108
rect 338724 3068 338730 3080
rect 339586 3068 339592 3080
rect 339644 3068 339650 3120
rect 347038 3068 347044 3120
rect 347096 3108 347102 3120
rect 354030 3108 354036 3120
rect 347096 3080 354036 3108
rect 347096 3068 347102 3080
rect 354030 3068 354036 3080
rect 354088 3068 354094 3120
rect 354140 3108 354168 3148
rect 354217 3145 354229 3179
rect 354263 3176 354275 3179
rect 355226 3176 355232 3188
rect 354263 3148 355232 3176
rect 354263 3145 354275 3148
rect 354217 3139 354275 3145
rect 355226 3136 355232 3148
rect 355284 3136 355290 3188
rect 364610 3176 364616 3188
rect 364306 3148 364616 3176
rect 357526 3108 357532 3120
rect 354140 3080 357532 3108
rect 357526 3068 357532 3080
rect 357584 3068 357590 3120
rect 358078 3068 358084 3120
rect 358136 3108 358142 3120
rect 363506 3108 363512 3120
rect 358136 3080 363512 3108
rect 358136 3068 358142 3080
rect 363506 3068 363512 3080
rect 363564 3068 363570 3120
rect 27706 3000 27712 3052
rect 27764 3040 27770 3052
rect 29638 3040 29644 3052
rect 27764 3012 29644 3040
rect 27764 3000 27770 3012
rect 29638 3000 29644 3012
rect 29696 3000 29702 3052
rect 103330 3000 103336 3052
rect 103388 3040 103394 3052
rect 266630 3040 266636 3052
rect 103388 3012 266636 3040
rect 103388 3000 103394 3012
rect 266630 3000 266636 3012
rect 266688 3000 266694 3052
rect 317322 3000 317328 3052
rect 317380 3040 317386 3052
rect 332962 3040 332968 3052
rect 317380 3012 332968 3040
rect 317380 3000 317386 3012
rect 332962 3000 332968 3012
rect 333020 3000 333026 3052
rect 348418 3000 348424 3052
rect 348476 3040 348482 3052
rect 354217 3043 354275 3049
rect 354217 3040 354229 3043
rect 348476 3012 354229 3040
rect 348476 3000 348482 3012
rect 354217 3009 354229 3012
rect 354263 3009 354275 3043
rect 354217 3003 354275 3009
rect 99834 2932 99840 2984
rect 99892 2972 99898 2984
rect 99892 2944 103514 2972
rect 99892 2932 99898 2944
rect 9950 2864 9956 2916
rect 10008 2904 10014 2916
rect 14458 2904 14464 2916
rect 10008 2876 14464 2904
rect 10008 2864 10014 2876
rect 14458 2864 14464 2876
rect 14516 2864 14522 2916
rect 103486 2904 103514 2944
rect 110506 2932 110512 2984
rect 110564 2972 110570 2984
rect 267918 2972 267924 2984
rect 110564 2944 267924 2972
rect 110564 2932 110570 2944
rect 267918 2932 267924 2944
rect 267976 2932 267982 2984
rect 304350 2932 304356 2984
rect 304408 2972 304414 2984
rect 304902 2972 304908 2984
rect 304408 2944 304908 2972
rect 304408 2932 304414 2944
rect 304902 2932 304908 2944
rect 304960 2932 304966 2984
rect 315022 2932 315028 2984
rect 315080 2972 315086 2984
rect 331674 2972 331680 2984
rect 315080 2944 331680 2972
rect 315080 2932 315086 2944
rect 331674 2932 331680 2944
rect 331732 2932 331738 2984
rect 336274 2932 336280 2984
rect 336332 2972 336338 2984
rect 338298 2972 338304 2984
rect 336332 2944 338304 2972
rect 336332 2932 336338 2944
rect 338298 2932 338304 2944
rect 338356 2932 338362 2984
rect 348510 2932 348516 2984
rect 348568 2972 348574 2984
rect 364306 2972 364334 3148
rect 364610 3136 364616 3148
rect 364668 3136 364674 3188
rect 375190 3136 375196 3188
rect 375248 3176 375254 3188
rect 454494 3176 454500 3188
rect 375248 3148 454500 3176
rect 375248 3136 375254 3148
rect 454494 3136 454500 3148
rect 454552 3136 454558 3188
rect 512638 3136 512644 3188
rect 512696 3176 512702 3188
rect 513558 3176 513564 3188
rect 512696 3148 513564 3176
rect 512696 3136 512702 3148
rect 513558 3136 513564 3148
rect 513616 3136 513622 3188
rect 373902 3068 373908 3120
rect 373960 3108 373966 3120
rect 447410 3108 447416 3120
rect 373960 3080 447416 3108
rect 373960 3068 373966 3080
rect 447410 3068 447416 3080
rect 447468 3068 447474 3120
rect 371142 3000 371148 3052
rect 371200 3040 371206 3052
rect 440234 3040 440240 3052
rect 371200 3012 440240 3040
rect 371200 3000 371206 3012
rect 440234 3000 440240 3012
rect 440292 3000 440298 3052
rect 440326 3000 440332 3052
rect 440384 3040 440390 3052
rect 441522 3040 441528 3052
rect 440384 3012 441528 3040
rect 440384 3000 440390 3012
rect 441522 3000 441528 3012
rect 441580 3000 441586 3052
rect 348568 2944 364334 2972
rect 348568 2932 348574 2944
rect 369762 2932 369768 2984
rect 369820 2972 369826 2984
rect 433242 2972 433248 2984
rect 369820 2944 433248 2972
rect 369820 2932 369826 2944
rect 433242 2932 433248 2944
rect 433300 2932 433306 2984
rect 111153 2907 111211 2913
rect 111153 2904 111165 2907
rect 103486 2876 111165 2904
rect 111153 2873 111165 2876
rect 111199 2873 111211 2907
rect 111153 2867 111211 2873
rect 114002 2864 114008 2916
rect 114060 2904 114066 2916
rect 114462 2904 114468 2916
rect 114060 2876 114468 2904
rect 114060 2864 114066 2876
rect 114462 2864 114468 2876
rect 114520 2864 114526 2916
rect 115198 2864 115204 2916
rect 115256 2904 115262 2916
rect 115842 2904 115848 2916
rect 115256 2876 115848 2904
rect 115256 2864 115262 2876
rect 115842 2864 115848 2876
rect 115900 2864 115906 2916
rect 116394 2864 116400 2916
rect 116452 2904 116458 2916
rect 117222 2904 117228 2916
rect 116452 2876 117228 2904
rect 116452 2864 116458 2876
rect 117222 2864 117228 2876
rect 117280 2864 117286 2916
rect 118786 2864 118792 2916
rect 118844 2904 118850 2916
rect 119798 2904 119804 2916
rect 118844 2876 119804 2904
rect 118844 2864 118850 2876
rect 119798 2864 119804 2876
rect 119856 2864 119862 2916
rect 122193 2907 122251 2913
rect 122193 2904 122205 2907
rect 119908 2876 122205 2904
rect 117590 2796 117596 2848
rect 117648 2836 117654 2848
rect 119908 2836 119936 2876
rect 122193 2873 122205 2876
rect 122239 2873 122251 2907
rect 122193 2867 122251 2873
rect 122282 2864 122288 2916
rect 122340 2904 122346 2916
rect 122742 2904 122748 2916
rect 122340 2876 122748 2904
rect 122340 2864 122346 2876
rect 122742 2864 122748 2876
rect 122800 2864 122806 2916
rect 123478 2864 123484 2916
rect 123536 2904 123542 2916
rect 124122 2904 124128 2916
rect 123536 2876 124128 2904
rect 123536 2864 123542 2876
rect 124122 2864 124128 2876
rect 124180 2864 124186 2916
rect 124674 2864 124680 2916
rect 124732 2904 124738 2916
rect 125410 2904 125416 2916
rect 124732 2876 125416 2904
rect 124732 2864 124738 2876
rect 125410 2864 125416 2876
rect 125468 2864 125474 2916
rect 270770 2904 270776 2916
rect 125612 2876 270776 2904
rect 117648 2808 119936 2836
rect 117648 2796 117654 2808
rect 121086 2796 121092 2848
rect 121144 2836 121150 2848
rect 125505 2839 125563 2845
rect 125505 2836 125517 2839
rect 121144 2808 122052 2836
rect 121144 2796 121150 2808
rect 122024 2700 122052 2808
rect 122300 2808 125517 2836
rect 122300 2700 122328 2808
rect 125505 2805 125517 2808
rect 125551 2805 125563 2839
rect 125505 2799 125563 2805
rect 122377 2771 122435 2777
rect 122377 2737 122389 2771
rect 122423 2768 122435 2771
rect 125612 2768 125640 2876
rect 270770 2864 270776 2876
rect 270828 2864 270834 2916
rect 316218 2864 316224 2916
rect 316276 2904 316282 2916
rect 331306 2904 331312 2916
rect 316276 2876 331312 2904
rect 316276 2864 316282 2876
rect 331306 2864 331312 2876
rect 331364 2864 331370 2916
rect 365622 2864 365628 2916
rect 365680 2904 365686 2916
rect 422570 2904 422576 2916
rect 365680 2876 422576 2904
rect 365680 2864 365686 2876
rect 422570 2864 422576 2876
rect 422628 2864 422634 2916
rect 125689 2839 125747 2845
rect 125689 2805 125701 2839
rect 125735 2836 125747 2839
rect 272058 2836 272064 2848
rect 125735 2808 272064 2836
rect 125735 2805 125747 2808
rect 125689 2799 125747 2805
rect 272058 2796 272064 2808
rect 272116 2796 272122 2848
rect 318518 2796 318524 2848
rect 318576 2836 318582 2848
rect 332778 2836 332784 2848
rect 318576 2808 332784 2836
rect 318576 2796 318582 2808
rect 332778 2796 332784 2808
rect 332836 2796 332842 2848
rect 364242 2796 364248 2848
rect 364300 2836 364306 2848
rect 415486 2836 415492 2848
rect 364300 2808 415492 2836
rect 364300 2796 364306 2808
rect 415486 2796 415492 2808
rect 415544 2796 415550 2848
rect 122423 2740 125640 2768
rect 122423 2737 122435 2740
rect 122377 2731 122435 2737
rect 122024 2672 122328 2700
rect 168374 1640 168380 1692
rect 168432 1680 168438 1692
rect 169662 1680 169668 1692
rect 168432 1652 169668 1680
rect 168432 1640 168438 1652
rect 169662 1640 169668 1652
rect 169720 1640 169726 1692
rect 456794 1368 456800 1420
rect 456852 1408 456858 1420
rect 458082 1408 458088 1420
rect 456852 1380 458088 1408
rect 456852 1368 456858 1380
rect 458082 1368 458088 1380
rect 458140 1368 458146 1420
<< via1 >>
rect 317328 700952 317380 701004
rect 429844 700952 429896 701004
rect 202788 700884 202840 700936
rect 331312 700884 331364 700936
rect 313188 700816 313240 700868
rect 462320 700816 462372 700868
rect 315948 700748 316000 700800
rect 478512 700748 478564 700800
rect 311808 700680 311860 700732
rect 494796 700680 494848 700732
rect 137836 700612 137888 700664
rect 336740 700612 336792 700664
rect 309048 700544 309100 700596
rect 527180 700544 527232 700596
rect 105452 700476 105504 700528
rect 106188 700476 106240 700528
rect 310428 700476 310480 700528
rect 543464 700476 543516 700528
rect 40500 700408 40552 700460
rect 41328 700408 41380 700460
rect 307668 700408 307720 700460
rect 559656 700408 559708 700460
rect 72976 700340 73028 700392
rect 340880 700340 340932 700392
rect 8116 700272 8168 700324
rect 345020 700272 345072 700324
rect 320088 700204 320140 700256
rect 413652 700204 413704 700256
rect 318708 700136 318760 700188
rect 397460 700136 397512 700188
rect 267648 700068 267700 700120
rect 327080 700068 327132 700120
rect 321468 700000 321520 700052
rect 364984 700000 365036 700052
rect 324228 699932 324280 699984
rect 348792 699932 348844 699984
rect 322848 699864 322900 699916
rect 332508 699864 332560 699916
rect 24308 699660 24360 699712
rect 24768 699660 24820 699712
rect 170312 699660 170364 699712
rect 171048 699660 171100 699712
rect 235172 699660 235224 699712
rect 235908 699660 235960 699712
rect 300124 699660 300176 699712
rect 300768 699660 300820 699712
rect 304908 696940 304960 696992
rect 580172 696940 580224 696992
rect 306288 683136 306340 683188
rect 580172 683136 580224 683188
rect 302148 670760 302200 670812
rect 580172 670760 580224 670812
rect 3516 670692 3568 670744
rect 333244 670692 333296 670744
rect 3516 656888 3568 656940
rect 350540 656888 350592 656940
rect 299388 643084 299440 643136
rect 580172 643084 580224 643136
rect 300676 630640 300728 630692
rect 580172 630640 580224 630692
rect 3332 618264 3384 618316
rect 338764 618264 338816 618316
rect 298008 616836 298060 616888
rect 580172 616836 580224 616888
rect 3332 605820 3384 605872
rect 354680 605820 354732 605872
rect 295248 590656 295300 590708
rect 579804 590656 579856 590708
rect 296628 576852 296680 576904
rect 580172 576852 580224 576904
rect 3056 565836 3108 565888
rect 342904 565836 342956 565888
rect 293868 563048 293920 563100
rect 579804 563048 579856 563100
rect 3332 553392 3384 553444
rect 360200 553392 360252 553444
rect 289728 536800 289780 536852
rect 580172 536800 580224 536852
rect 291108 524424 291160 524476
rect 580172 524424 580224 524476
rect 3332 514768 3384 514820
rect 348424 514768 348476 514820
rect 288348 510620 288400 510672
rect 580172 510620 580224 510672
rect 3240 500964 3292 501016
rect 364340 500964 364392 501016
rect 285588 484372 285640 484424
rect 580172 484372 580224 484424
rect 286968 470568 287020 470620
rect 579988 470568 580040 470620
rect 3516 462340 3568 462392
rect 352564 462340 352616 462392
rect 171048 460844 171100 460896
rect 334900 460844 334952 460896
rect 154488 460776 154540 460828
rect 338120 460776 338172 460828
rect 338764 460776 338816 460828
rect 356980 460776 357032 460828
rect 106188 460708 106240 460760
rect 339684 460708 339736 460760
rect 89628 460640 89680 460692
rect 342812 460640 342864 460692
rect 342904 460640 342956 460692
rect 361764 460640 361816 460692
rect 41328 460572 41380 460624
rect 344376 460572 344428 460624
rect 24768 460504 24820 460556
rect 347780 460504 347832 460556
rect 348424 460504 348476 460556
rect 366456 460504 366508 460556
rect 3424 460436 3476 460488
rect 349160 460436 349212 460488
rect 352564 460436 352616 460488
rect 371240 460436 371292 460488
rect 3608 460368 3660 460420
rect 353852 460368 353904 460420
rect 3700 460300 3752 460352
rect 358820 460300 358872 460352
rect 3792 460232 3844 460284
rect 363328 460232 363380 460284
rect 3884 460164 3936 460216
rect 368112 460164 368164 460216
rect 219348 460096 219400 460148
rect 235908 460028 235960 460080
rect 330208 460028 330260 460080
rect 333244 460096 333296 460148
rect 352288 460096 352340 460148
rect 333336 460028 333388 460080
rect 284208 459960 284260 460012
rect 328552 459960 328604 460012
rect 300768 459824 300820 459876
rect 325700 459892 325752 459944
rect 281448 459756 281500 459808
rect 285036 459688 285088 459740
rect 285588 459688 285640 459740
rect 292948 459756 293000 459808
rect 293868 459756 293920 459808
rect 294512 459756 294564 459808
rect 295248 459756 295300 459808
rect 296076 459756 296128 459808
rect 296628 459756 296680 459808
rect 303988 459756 304040 459808
rect 304908 459756 304960 459808
rect 305552 459756 305604 459808
rect 306288 459756 306340 459808
rect 307116 459756 307168 459808
rect 307668 459756 307720 459808
rect 315028 459756 315080 459808
rect 315948 459756 316000 459808
rect 316592 459756 316644 459808
rect 317328 459756 317380 459808
rect 318156 459756 318208 459808
rect 318708 459756 318760 459808
rect 569224 459688 569276 459740
rect 272340 459620 272392 459672
rect 566464 459620 566516 459672
rect 267464 459552 267516 459604
rect 562324 459552 562376 459604
rect 273996 458804 274048 458856
rect 416044 458804 416096 458856
rect 231124 458736 231176 458788
rect 374368 458736 374420 458788
rect 280068 458668 280120 458720
rect 429844 458668 429896 458720
rect 222844 458600 222896 458652
rect 375932 458600 375984 458652
rect 277032 458532 277084 458584
rect 432604 458532 432656 458584
rect 232596 458464 232648 458516
rect 391940 458464 391992 458516
rect 270408 458396 270460 458448
rect 428556 458396 428608 458448
rect 228364 458328 228416 458380
rect 407580 458328 407632 458380
rect 269028 458260 269080 458312
rect 580264 458260 580316 458312
rect 3424 458192 3476 458244
rect 373126 458192 373178 458244
rect 283472 457487 283524 457496
rect 283472 457453 283481 457487
rect 283481 457453 283515 457487
rect 283515 457453 283524 457487
rect 283472 457444 283524 457453
rect 233884 457376 233936 457428
rect 369860 457376 369912 457428
rect 377588 457419 377640 457428
rect 377588 457385 377597 457419
rect 377597 457385 377631 457419
rect 377631 457385 377640 457419
rect 377588 457376 377640 457385
rect 379152 457419 379204 457428
rect 379152 457385 379161 457419
rect 379161 457385 379195 457419
rect 379195 457385 379204 457419
rect 379152 457376 379204 457385
rect 380900 457419 380952 457428
rect 380900 457385 380909 457419
rect 380909 457385 380943 457419
rect 380943 457385 380952 457419
rect 380900 457376 380952 457385
rect 278688 457308 278740 457360
rect 418804 457308 418856 457360
rect 239220 457283 239272 457292
rect 239220 457249 239229 457283
rect 239229 457249 239263 457283
rect 239263 457249 239272 457283
rect 239220 457240 239272 457249
rect 255044 457283 255096 457292
rect 255044 457249 255053 457283
rect 255053 457249 255087 457283
rect 255087 457249 255096 457283
rect 255044 457240 255096 457249
rect 266084 457283 266136 457292
rect 266084 457249 266093 457283
rect 266093 457249 266127 457283
rect 266127 457249 266136 457283
rect 266084 457240 266136 457249
rect 275560 457240 275612 457292
rect 425704 457240 425756 457292
rect 226984 457172 227036 457224
rect 421656 457104 421708 457156
rect 224224 457036 224276 457088
rect 417424 456968 417476 457020
rect 431224 456900 431276 456952
rect 579804 456832 579856 456884
rect 4804 456764 4856 456816
rect 3332 449828 3384 449880
rect 233884 449828 233936 449880
rect 429844 431876 429896 431928
rect 580172 431876 580224 431928
rect 569224 419432 569276 419484
rect 580172 419432 580224 419484
rect 3424 411204 3476 411256
rect 222844 411204 222896 411256
rect 418804 405628 418856 405680
rect 579620 405628 579672 405680
rect 3240 398760 3292 398812
rect 231124 398760 231176 398812
rect 425704 379448 425756 379500
rect 580172 379448 580224 379500
rect 2780 371424 2832 371476
rect 4804 371424 4856 371476
rect 432604 365644 432656 365696
rect 580172 365644 580224 365696
rect 3332 358708 3384 358760
rect 224224 358708 224276 358760
rect 416044 353200 416096 353252
rect 580172 353200 580224 353252
rect 3148 346332 3200 346384
rect 226984 346332 227036 346384
rect 220084 336676 220136 336728
rect 288532 336676 288584 336728
rect 289820 336676 289872 336728
rect 310520 336744 310572 336796
rect 310796 336744 310848 336796
rect 215944 336608 215996 336660
rect 214564 336540 214616 336592
rect 288440 336608 288492 336660
rect 290004 336608 290056 336660
rect 291384 336676 291436 336728
rect 292948 336676 293000 336728
rect 300492 336676 300544 336728
rect 301320 336676 301372 336728
rect 304908 336676 304960 336728
rect 328736 336676 328788 336728
rect 329196 336676 329248 336728
rect 333980 336676 334032 336728
rect 339500 336676 339552 336728
rect 339776 336676 339828 336728
rect 341616 336676 341668 336728
rect 342076 336676 342128 336728
rect 343548 336676 343600 336728
rect 344284 336676 344336 336728
rect 347044 336676 347096 336728
rect 347688 336676 347740 336728
rect 348148 336676 348200 336728
rect 349068 336676 349120 336728
rect 351092 336676 351144 336728
rect 351828 336676 351880 336728
rect 352840 336676 352892 336728
rect 353116 336676 353168 336728
rect 355692 336676 355744 336728
rect 355968 336676 356020 336728
rect 357164 336676 357216 336728
rect 357348 336676 357400 336728
rect 358360 336676 358412 336728
rect 358636 336676 358688 336728
rect 360568 336676 360620 336728
rect 361120 336676 361172 336728
rect 362592 336676 362644 336728
rect 362868 336676 362920 336728
rect 363512 336676 363564 336728
rect 364248 336676 364300 336728
rect 367468 336676 367520 336728
rect 368296 336676 368348 336728
rect 368940 336676 368992 336728
rect 369768 336676 369820 336728
rect 369860 336676 369912 336728
rect 436100 336676 436152 336728
rect 294420 336608 294472 336660
rect 296536 336608 296588 336660
rect 296904 336608 296956 336660
rect 300768 336608 300820 336660
rect 327540 336608 327592 336660
rect 355048 336608 355100 336660
rect 355876 336608 355928 336660
rect 292212 336540 292264 336592
rect 296628 336540 296680 336592
rect 326160 336540 326212 336592
rect 327724 336540 327776 336592
rect 328460 336540 328512 336592
rect 348424 336540 348476 336592
rect 356888 336540 356940 336592
rect 357348 336540 357400 336592
rect 357992 336608 358044 336660
rect 358728 336608 358780 336660
rect 362040 336608 362092 336660
rect 362684 336608 362736 336660
rect 366456 336608 366508 336660
rect 367008 336608 367060 336660
rect 372252 336608 372304 336660
rect 443000 336608 443052 336660
rect 363604 336540 363656 336592
rect 373356 336540 373408 336592
rect 373908 336540 373960 336592
rect 375932 336540 375984 336592
rect 376668 336540 376720 336592
rect 377036 336540 377088 336592
rect 377864 336540 377916 336592
rect 380256 336540 380308 336592
rect 380716 336540 380768 336592
rect 382004 336540 382056 336592
rect 382188 336540 382240 336592
rect 449900 336540 449952 336592
rect 209044 336472 209096 336524
rect 296720 336472 296772 336524
rect 299388 336472 299440 336524
rect 327080 336472 327132 336524
rect 347412 336472 347464 336524
rect 358084 336472 358136 336524
rect 367836 336472 367888 336524
rect 379888 336472 379940 336524
rect 380808 336472 380860 336524
rect 381360 336472 381412 336524
rect 381912 336472 381964 336524
rect 125508 336404 125560 336456
rect 273260 336404 273312 336456
rect 276020 336404 276072 336456
rect 279056 336404 279108 336456
rect 282644 336404 282696 336456
rect 283380 336404 283432 336456
rect 293316 336404 293368 336456
rect 323584 336404 323636 336456
rect 352196 336404 352248 336456
rect 369308 336404 369360 336456
rect 456800 336472 456852 336524
rect 114468 336336 114520 336388
rect 269948 336336 270000 336388
rect 277308 336336 277360 336388
rect 319904 336336 319956 336388
rect 346676 336336 346728 336388
rect 347596 336336 347648 336388
rect 354404 336336 354456 336388
rect 370504 336336 370556 336388
rect 376576 336336 376628 336388
rect 383936 336404 383988 336456
rect 384856 336404 384908 336456
rect 387248 336404 387300 336456
rect 387708 336404 387760 336456
rect 388352 336404 388404 336456
rect 389088 336404 389140 336456
rect 389456 336404 389508 336456
rect 390192 336404 390244 336456
rect 392676 336404 392728 336456
rect 393136 336404 393188 336456
rect 465080 336404 465132 336456
rect 381728 336336 381780 336388
rect 468484 336336 468536 336388
rect 107568 336268 107620 336320
rect 267832 336268 267884 336320
rect 277400 336268 277452 336320
rect 279792 336268 279844 336320
rect 282184 336268 282236 336320
rect 283104 336268 283156 336320
rect 321560 336268 321612 336320
rect 346308 336268 346360 336320
rect 347136 336268 347188 336320
rect 348884 336268 348936 336320
rect 367468 336268 367520 336320
rect 380992 336268 381044 336320
rect 471980 336268 472032 336320
rect 57244 336200 57296 336252
rect 251272 336200 251324 336252
rect 259460 336200 259512 336252
rect 261484 336200 261536 336252
rect 264520 336200 264572 336252
rect 265164 336200 265216 336252
rect 270040 336200 270092 336252
rect 271880 336200 271932 336252
rect 274548 336200 274600 336252
rect 319260 336200 319312 336252
rect 354036 336200 354088 336252
rect 354496 336200 354548 336252
rect 371792 336200 371844 336252
rect 374460 336200 374512 336252
rect 383476 336200 383528 336252
rect 475384 336200 475436 336252
rect 51724 336132 51776 336184
rect 247960 336132 248012 336184
rect 267648 336132 267700 336184
rect 317052 336132 317104 336184
rect 344100 336132 344152 336184
rect 345664 336132 345716 336184
rect 351460 336132 351512 336184
rect 375472 336132 375524 336184
rect 50344 336064 50396 336116
rect 245844 336064 245896 336116
rect 270408 336064 270460 336116
rect 318156 336064 318208 336116
rect 328368 336064 328420 336116
rect 336004 336064 336056 336116
rect 353668 336064 353720 336116
rect 382464 336132 382516 336184
rect 383200 336132 383252 336184
rect 478880 336132 478932 336184
rect 378876 336064 378928 336116
rect 393228 336064 393280 336116
rect 497464 336064 497516 336116
rect 35164 335996 35216 336048
rect 243636 335996 243688 336048
rect 263508 335996 263560 336048
rect 316040 335996 316092 336048
rect 316684 335996 316736 336048
rect 327264 335996 327316 336048
rect 333244 335996 333296 336048
rect 336740 335996 336792 336048
rect 344836 335996 344888 336048
rect 348424 335996 348476 336048
rect 356520 335996 356572 336048
rect 388444 335996 388496 336048
rect 391204 335996 391256 336048
rect 504364 335996 504416 336048
rect 204904 335928 204956 335980
rect 276848 335928 276900 335980
rect 281356 335928 281408 335980
rect 286416 335928 286468 335980
rect 315212 335928 315264 335980
rect 336004 335928 336056 335980
rect 337476 335928 337528 335980
rect 370412 335928 370464 335980
rect 435364 335928 435416 335980
rect 224224 335860 224276 335912
rect 291200 335860 291252 335912
rect 291936 335860 291988 335912
rect 311900 335860 311952 335912
rect 366916 335860 366968 335912
rect 233884 335792 233936 335844
rect 300216 335792 300268 335844
rect 345572 335792 345624 335844
rect 349804 335792 349856 335844
rect 359096 335792 359148 335844
rect 360016 335792 360068 335844
rect 371884 335792 371936 335844
rect 372344 335792 372396 335844
rect 372988 335860 373040 335912
rect 374644 335860 374696 335912
rect 429200 335860 429252 335912
rect 425704 335792 425756 335844
rect 222844 335724 222896 335776
rect 287796 335724 287848 335776
rect 289084 335724 289136 335776
rect 313004 335724 313056 335776
rect 352564 335724 352616 335776
rect 353208 335724 353260 335776
rect 428464 335724 428516 335776
rect 226984 335656 227036 335708
rect 288900 335656 288952 335708
rect 295984 335656 296036 335708
rect 314936 335656 314988 335708
rect 342720 335656 342772 335708
rect 343364 335656 343416 335708
rect 349620 335656 349672 335708
rect 353944 335656 353996 335708
rect 361212 335656 361264 335708
rect 361488 335656 361540 335708
rect 366824 335656 366876 335708
rect 425060 335656 425112 335708
rect 213184 335588 213236 335640
rect 273904 335588 273956 335640
rect 288348 335588 288400 335640
rect 296444 335588 296496 335640
rect 298100 335588 298152 335640
rect 366088 335588 366140 335640
rect 413192 335588 413244 335640
rect 413836 335588 413888 335640
rect 414848 335588 414900 335640
rect 415124 335588 415176 335640
rect 421564 335588 421616 335640
rect 231124 335520 231176 335572
rect 285680 335520 285732 335572
rect 341248 335520 341300 335572
rect 342352 335520 342404 335572
rect 347504 335520 347556 335572
rect 348516 335520 348568 335572
rect 364984 335520 365036 335572
rect 414664 335520 414716 335572
rect 415308 335520 415360 335572
rect 232504 335452 232556 335504
rect 282368 335452 282420 335504
rect 344468 335452 344520 335504
rect 346952 335452 347004 335504
rect 363880 335452 363932 335504
rect 416780 335452 416832 335504
rect 233976 335384 234028 335436
rect 273536 335384 273588 335436
rect 341984 335384 342036 335436
rect 345112 335384 345164 335436
rect 350080 335384 350132 335436
rect 350356 335384 350408 335436
rect 364616 335384 364668 335436
rect 418160 335384 418212 335436
rect 267740 335316 267792 335368
rect 272800 335316 272852 335368
rect 274456 335316 274508 335368
rect 278780 335316 278832 335368
rect 197268 335248 197320 335300
rect 295432 335316 295484 335368
rect 332508 335316 332560 335368
rect 337108 335316 337160 335368
rect 344928 335316 344980 335368
rect 345756 335316 345808 335368
rect 355416 335316 355468 335368
rect 382924 335316 382976 335368
rect 384672 335316 384724 335368
rect 388996 335316 389048 335368
rect 393228 335316 393280 335368
rect 397828 335316 397880 335368
rect 398564 335316 398616 335368
rect 402244 335316 402296 335368
rect 402704 335316 402756 335368
rect 403992 335316 404044 335368
rect 404268 335316 404320 335368
rect 405188 335316 405240 335368
rect 405556 335316 405608 335368
rect 406568 335316 406620 335368
rect 406844 335316 406896 335368
rect 407672 335316 407724 335368
rect 408316 335316 408368 335368
rect 409512 335316 409564 335368
rect 409788 335316 409840 335368
rect 410708 335316 410760 335368
rect 411076 335316 411128 335368
rect 412088 335316 412140 335368
rect 412364 335316 412416 335368
rect 418804 335316 418856 335368
rect 373724 335248 373776 335300
rect 448520 335248 448572 335300
rect 179328 335180 179380 335232
rect 288440 335180 288492 335232
rect 483020 335180 483072 335232
rect 169668 335112 169720 335164
rect 286692 335112 286744 335164
rect 384304 335112 384356 335164
rect 481640 335112 481692 335164
rect 161388 335044 161440 335096
rect 284484 335044 284536 335096
rect 391940 335044 391992 335096
rect 490012 335044 490064 335096
rect 144828 334976 144880 335028
rect 276020 334976 276072 335028
rect 390100 334976 390152 335028
rect 500960 334976 501012 335028
rect 147588 334908 147640 334960
rect 280252 334908 280304 334960
rect 392308 334908 392360 334960
rect 507860 334908 507912 334960
rect 140688 334840 140740 334892
rect 277952 334840 278004 334892
rect 393780 334840 393832 334892
rect 512644 334840 512696 334892
rect 87604 334772 87656 334824
rect 260932 334772 260984 334824
rect 398196 334772 398248 334824
rect 526444 334772 526496 334824
rect 86868 334704 86920 334756
rect 259460 334704 259512 334756
rect 397092 334704 397144 334756
rect 522304 334704 522356 334756
rect 29644 334636 29696 334688
rect 243268 334636 243320 334688
rect 398472 334636 398524 334688
rect 528560 334636 528612 334688
rect 22744 334568 22796 334620
rect 238852 334568 238904 334620
rect 402520 334568 402572 334620
rect 540244 334568 540296 334620
rect 202788 334500 202840 334552
rect 296536 334500 296588 334552
rect 371516 334500 371568 334552
rect 440332 334500 440384 334552
rect 216588 334432 216640 334484
rect 300492 334432 300544 334484
rect 368112 334432 368164 334484
rect 430580 334432 430632 334484
rect 223488 334364 223540 334416
rect 303620 334364 303672 334416
rect 205548 333888 205600 333940
rect 296444 333888 296496 333940
rect 374644 333888 374696 333940
rect 445760 333888 445812 333940
rect 198648 333820 198700 333872
rect 295800 333820 295852 333872
rect 373816 333820 373868 333872
rect 448612 333820 448664 333872
rect 177948 333752 178000 333804
rect 288532 333752 288584 333804
rect 377404 333752 377456 333804
rect 459560 333752 459612 333804
rect 162768 333684 162820 333736
rect 284852 333684 284904 333736
rect 380900 333684 380952 333736
rect 470600 333684 470652 333736
rect 158628 333616 158680 333668
rect 282644 333616 282696 333668
rect 387616 333616 387668 333668
rect 492680 333616 492732 333668
rect 151728 333548 151780 333600
rect 281448 333548 281500 333600
rect 390928 333548 390980 333600
rect 502984 333548 503036 333600
rect 93124 333480 93176 333532
rect 262956 333480 263008 333532
rect 394608 333480 394660 333532
rect 515404 333480 515456 333532
rect 88984 333412 89036 333464
rect 261944 333412 261996 333464
rect 395896 333412 395948 333464
rect 520280 333412 520332 333464
rect 84108 333344 84160 333396
rect 260380 333344 260432 333396
rect 400128 333344 400180 333396
rect 54484 333276 54536 333328
rect 247592 333276 247644 333328
rect 530584 333344 530636 333396
rect 533344 333276 533396 333328
rect 39304 333208 39356 333260
rect 241888 333208 241940 333260
rect 401508 333208 401560 333260
rect 538220 333208 538272 333260
rect 209688 333140 209740 333192
rect 299112 333140 299164 333192
rect 399300 333140 399352 333192
rect 227628 333072 227680 333124
rect 304632 333072 304684 333124
rect 219256 332528 219308 332580
rect 302424 332528 302476 332580
rect 188988 332460 189040 332512
rect 291384 332460 291436 332512
rect 182088 332392 182140 332444
rect 290832 332392 290884 332444
rect 375196 332392 375248 332444
rect 452660 332392 452712 332444
rect 175188 332324 175240 332376
rect 288624 332324 288676 332376
rect 376208 332324 376260 332376
rect 456892 332324 456944 332376
rect 171048 332256 171100 332308
rect 287428 332256 287480 332308
rect 378508 332256 378560 332308
rect 463700 332256 463752 332308
rect 143448 332188 143500 332240
rect 274456 332188 274508 332240
rect 379428 332188 379480 332240
rect 466460 332188 466512 332240
rect 104164 332120 104216 332172
rect 266360 332120 266412 332172
rect 382832 332120 382884 332172
rect 477500 332120 477552 332172
rect 99288 332052 99340 332104
rect 264520 332052 264572 332104
rect 385316 332052 385368 332104
rect 485780 332052 485832 332104
rect 95148 331984 95200 332036
rect 264060 331984 264112 332036
rect 388720 331984 388772 332036
rect 496820 331984 496872 332036
rect 68284 331916 68336 331968
rect 250168 331916 250220 331968
rect 391848 331916 391900 331968
rect 506480 331916 506532 331968
rect 33784 331848 33836 331900
rect 244464 331848 244516 331900
rect 396356 331848 396408 331900
rect 519544 331848 519596 331900
rect 153108 330964 153160 331016
rect 282000 330964 282052 331016
rect 146208 330896 146260 330948
rect 277400 330896 277452 330948
rect 117228 330828 117280 330880
rect 270868 330828 270920 330880
rect 399668 330828 399720 330880
rect 485044 330828 485096 330880
rect 111064 330760 111116 330812
rect 268476 330760 268528 330812
rect 324412 330760 324464 330812
rect 386328 330760 386380 330812
rect 489184 330760 489236 330812
rect 106188 330692 106240 330744
rect 267372 330692 267424 330744
rect 81348 330624 81400 330676
rect 259644 330624 259696 330676
rect 389824 330692 389876 330744
rect 499580 330692 499632 330744
rect 392860 330624 392912 330676
rect 510620 330624 510672 330676
rect 58624 330556 58676 330608
rect 248696 330556 248748 330608
rect 324412 330556 324464 330608
rect 394148 330556 394200 330608
rect 514760 330556 514812 330608
rect 36544 330488 36596 330540
rect 234804 330420 234856 330472
rect 235540 330420 235592 330472
rect 236092 330420 236144 330472
rect 237012 330420 237064 330472
rect 237380 330420 237432 330472
rect 238484 330420 238536 330472
rect 241612 330488 241664 330540
rect 242532 330488 242584 330540
rect 244372 330488 244424 330540
rect 245108 330488 245160 330540
rect 247132 330488 247184 330540
rect 247316 330488 247368 330540
rect 248512 330488 248564 330540
rect 249432 330488 249484 330540
rect 249892 330488 249944 330540
rect 250904 330488 250956 330540
rect 251272 330488 251324 330540
rect 252008 330488 252060 330540
rect 253940 330488 253992 330540
rect 254584 330488 254636 330540
rect 255412 330488 255464 330540
rect 256056 330488 256108 330540
rect 258172 330488 258224 330540
rect 259000 330488 259052 330540
rect 262404 330488 262456 330540
rect 262588 330488 262640 330540
rect 265164 330488 265216 330540
rect 265900 330488 265952 330540
rect 266452 330488 266504 330540
rect 267004 330488 267056 330540
rect 270592 330488 270644 330540
rect 271328 330488 271380 330540
rect 285772 330488 285824 330540
rect 286324 330488 286376 330540
rect 287152 330488 287204 330540
rect 288164 330488 288216 330540
rect 291292 330488 291344 330540
rect 291844 330488 291896 330540
rect 294052 330488 294104 330540
rect 295156 330488 295208 330540
rect 300952 330488 301004 330540
rect 301688 330488 301740 330540
rect 305092 330488 305144 330540
rect 305736 330488 305788 330540
rect 307760 330488 307812 330540
rect 308588 330488 308640 330540
rect 309324 330488 309376 330540
rect 310060 330488 310112 330540
rect 310612 330488 310664 330540
rect 311164 330488 311216 330540
rect 311992 330488 312044 330540
rect 312636 330488 312688 330540
rect 313280 330488 313332 330540
rect 314108 330488 314160 330540
rect 317604 330488 317656 330540
rect 318524 330488 318576 330540
rect 318892 330488 318944 330540
rect 319536 330488 319588 330540
rect 320272 330488 320324 330540
rect 321008 330488 321060 330540
rect 321652 330488 321704 330540
rect 322112 330488 322164 330540
rect 323124 330488 323176 330540
rect 323952 330488 324004 330540
rect 324504 330488 324556 330540
rect 325424 330488 325476 330540
rect 325792 330488 325844 330540
rect 326528 330488 326580 330540
rect 328552 330488 328604 330540
rect 329472 330488 329524 330540
rect 330024 330488 330076 330540
rect 330576 330488 330628 330540
rect 331312 330488 331364 330540
rect 332324 330488 332376 330540
rect 332692 330488 332744 330540
rect 333428 330488 333480 330540
rect 334072 330488 334124 330540
rect 334532 330488 334584 330540
rect 335544 330488 335596 330540
rect 336372 330488 336424 330540
rect 338120 330488 338172 330540
rect 338948 330488 339000 330540
rect 349988 330488 350040 330540
rect 350448 330488 350500 330540
rect 401876 330488 401928 330540
rect 402796 330488 402848 330540
rect 245660 330420 245712 330472
rect 254032 330420 254084 330472
rect 254952 330420 255004 330472
rect 262312 330420 262364 330472
rect 263324 330420 263376 330472
rect 305184 330420 305236 330472
rect 306104 330420 306156 330472
rect 309140 330420 309192 330472
rect 309692 330420 309744 330472
rect 329932 330420 329984 330472
rect 330944 330420 330996 330472
rect 395252 330420 395304 330472
rect 517520 330488 517572 330540
rect 403256 330420 403308 330472
rect 404176 330420 404228 330472
rect 404728 330420 404780 330472
rect 405464 330420 405516 330472
rect 406200 330420 406252 330472
rect 406936 330420 406988 330472
rect 408776 330420 408828 330472
rect 409696 330420 409748 330472
rect 410248 330420 410300 330472
rect 410984 330420 411036 330472
rect 411720 330420 411772 330472
rect 412548 330420 412600 330472
rect 414296 330420 414348 330472
rect 415216 330420 415268 330472
rect 405096 330352 405148 330404
rect 405648 330352 405700 330404
rect 410616 330352 410668 330404
rect 411168 330352 411220 330404
rect 332600 330148 332652 330200
rect 333060 330148 333112 330200
rect 299572 330012 299624 330064
rect 300584 330012 300636 330064
rect 271972 329808 272024 329860
rect 272432 329808 272484 329860
rect 255320 329604 255372 329656
rect 255688 329604 255740 329656
rect 124128 329400 124180 329452
rect 267740 329400 267792 329452
rect 119988 329332 120040 329384
rect 270040 329332 270092 329384
rect 113088 329264 113140 329316
rect 269580 329264 269632 329316
rect 61384 329196 61436 329248
rect 252560 329196 252612 329248
rect 47584 329128 47636 329180
rect 246580 329128 246632 329180
rect 397368 329128 397420 329180
rect 524420 329128 524472 329180
rect 32404 329060 32456 329112
rect 240324 329060 240376 329112
rect 400772 329060 400824 329112
rect 535460 329060 535512 329112
rect 14464 327700 14516 327752
rect 237748 327700 237800 327752
rect 314752 327156 314804 327208
rect 315580 327156 315632 327208
rect 305000 326884 305052 326936
rect 305368 326884 305420 326936
rect 334164 326680 334216 326732
rect 334900 326680 334952 326732
rect 306472 326476 306524 326528
rect 307484 326476 307536 326528
rect 276204 326408 276256 326460
rect 274640 326340 274692 326392
rect 275744 326340 275796 326392
rect 277492 326340 277544 326392
rect 277676 326340 277728 326392
rect 280252 326340 280304 326392
rect 280896 326340 280948 326392
rect 360936 326340 360988 326392
rect 361304 326340 361356 326392
rect 362408 326340 362460 326392
rect 362868 326340 362920 326392
rect 276204 326204 276256 326256
rect 428556 325592 428608 325644
rect 579896 325592 579948 325644
rect 277492 325116 277544 325168
rect 278320 325116 278372 325168
rect 276112 323620 276164 323672
rect 276296 323620 276348 323672
rect 566464 313216 566516 313268
rect 580172 313216 580224 313268
rect 421656 273164 421708 273216
rect 580172 273164 580224 273216
rect 562324 259360 562376 259412
rect 580172 259360 580224 259412
rect 3332 215228 3384 215280
rect 232596 215228 232648 215280
rect 417424 166948 417476 167000
rect 580172 166948 580224 167000
rect 3424 45500 3476 45552
rect 228364 45500 228416 45552
rect 3424 20612 3476 20664
rect 414940 20612 414992 20664
rect 431224 20612 431276 20664
rect 579988 20612 580040 20664
rect 157248 18572 157300 18624
rect 282184 18572 282236 18624
rect 161296 17212 161348 17264
rect 284392 17212 284444 17264
rect 138848 15852 138900 15904
rect 277584 15852 277636 15904
rect 252376 14424 252428 14476
rect 311992 14424 312044 14476
rect 186136 13336 186188 13388
rect 291292 13336 291344 13388
rect 125876 13268 125928 13320
rect 233976 13268 234028 13320
rect 163688 13200 163740 13252
rect 284484 13200 284536 13252
rect 149520 13132 149572 13184
rect 280252 13132 280304 13184
rect 128176 13064 128228 13116
rect 273444 13064 273496 13116
rect 212172 12180 212224 12232
rect 233884 12180 233936 12232
rect 182548 12112 182600 12164
rect 224224 12112 224276 12164
rect 175464 12044 175516 12096
rect 226984 12044 227036 12096
rect 164884 11976 164936 12028
rect 231124 11976 231176 12028
rect 154212 11908 154264 11960
rect 232504 11908 232556 11960
rect 251088 11908 251140 11960
rect 291844 11908 291896 11960
rect 167184 11840 167236 11892
rect 285772 11840 285824 11892
rect 78588 11772 78640 11824
rect 258356 11772 258408 11824
rect 74448 11704 74500 11756
rect 256884 11704 256936 11756
rect 448612 11704 448664 11756
rect 449808 11704 449860 11756
rect 160100 11636 160152 11688
rect 161296 11636 161348 11688
rect 95056 10956 95108 11008
rect 263692 10956 263744 11008
rect 91008 10888 91060 10940
rect 262404 10888 262456 10940
rect 70308 10820 70360 10872
rect 255596 10820 255648 10872
rect 67548 10752 67600 10804
rect 255504 10752 255556 10804
rect 63224 10684 63276 10736
rect 254216 10684 254268 10736
rect 60648 10616 60700 10668
rect 252744 10616 252796 10668
rect 260656 10616 260708 10668
rect 286324 10616 286376 10668
rect 56508 10548 56560 10600
rect 251272 10548 251324 10600
rect 253480 10548 253532 10600
rect 289084 10548 289136 10600
rect 53748 10480 53800 10532
rect 249892 10480 249944 10532
rect 271788 10480 271840 10532
rect 317604 10480 317656 10532
rect 49608 10412 49660 10464
rect 249984 10412 250036 10464
rect 269028 10412 269080 10464
rect 317512 10412 317564 10464
rect 45468 10344 45520 10396
rect 248604 10344 248656 10396
rect 264888 10344 264940 10396
rect 316132 10344 316184 10396
rect 41328 10276 41380 10328
rect 247132 10276 247184 10328
rect 256608 10276 256660 10328
rect 313464 10276 313516 10328
rect 353024 10276 353076 10328
rect 382372 10276 382424 10328
rect 382924 10276 382976 10328
rect 389456 10276 389508 10328
rect 97908 10208 97960 10260
rect 265072 10208 265124 10260
rect 102048 10140 102100 10192
rect 265164 10140 265216 10192
rect 104532 10072 104584 10124
rect 266452 10072 266504 10124
rect 108948 10004 109000 10056
rect 267832 10004 267884 10056
rect 111616 9936 111668 9988
rect 269304 9936 269356 9988
rect 115848 9868 115900 9920
rect 270684 9868 270736 9920
rect 119804 9800 119856 9852
rect 270592 9800 270644 9852
rect 122748 9732 122800 9784
rect 271972 9732 272024 9784
rect 209780 9596 209832 9648
rect 299664 9596 299716 9648
rect 206192 9528 206244 9580
rect 298192 9528 298244 9580
rect 202696 9460 202748 9512
rect 296812 9460 296864 9512
rect 199108 9392 199160 9444
rect 295524 9392 295576 9444
rect 195612 9324 195664 9376
rect 294052 9324 294104 9376
rect 192024 9256 192076 9308
rect 294144 9256 294196 9308
rect 135260 9188 135312 9240
rect 276112 9188 276164 9240
rect 131764 9120 131816 9172
rect 274916 9120 274968 9172
rect 37188 9052 37240 9104
rect 245844 9052 245896 9104
rect 248788 9052 248840 9104
rect 310796 9052 310848 9104
rect 33600 8984 33652 9036
rect 244372 8984 244424 9036
rect 245200 8984 245252 9036
rect 310704 8984 310756 9036
rect 357164 8984 357216 9036
rect 396540 8984 396592 9036
rect 432604 8984 432656 9036
rect 494704 8984 494756 9036
rect 8760 8916 8812 8968
rect 237472 8916 237524 8968
rect 238116 8916 238168 8968
rect 307944 8916 307996 8968
rect 353944 8916 353996 8968
rect 370596 8916 370648 8968
rect 372436 8916 372488 8968
rect 445024 8916 445076 8968
rect 126980 8848 127032 8900
rect 213184 8848 213236 8900
rect 213368 8848 213420 8900
rect 299572 8848 299624 8900
rect 216864 8780 216916 8832
rect 300952 8780 301004 8832
rect 220452 8712 220504 8764
rect 302424 8712 302476 8764
rect 223948 8644 224000 8696
rect 303712 8644 303764 8696
rect 227536 8576 227588 8628
rect 305276 8576 305328 8628
rect 231032 8508 231084 8560
rect 305184 8508 305236 8560
rect 234988 8440 235040 8492
rect 306656 8440 306708 8492
rect 241704 8372 241756 8424
rect 309416 8372 309468 8424
rect 421564 8304 421616 8356
rect 423772 8304 423824 8356
rect 428464 8304 428516 8356
rect 434444 8304 434496 8356
rect 137652 8236 137704 8288
rect 277676 8236 277728 8288
rect 372344 8236 372396 8288
rect 442632 8236 442684 8288
rect 134156 8168 134208 8220
rect 276204 8168 276256 8220
rect 403992 8168 404044 8220
rect 545488 8168 545540 8220
rect 79692 8100 79744 8152
rect 76196 8032 76248 8084
rect 258356 8100 258408 8152
rect 259552 8100 259604 8152
rect 265348 8100 265400 8152
rect 316224 8100 316276 8152
rect 405464 8100 405516 8152
rect 549076 8100 549128 8152
rect 258264 8032 258316 8084
rect 72608 7964 72660 8016
rect 256792 7964 256844 8016
rect 261760 8032 261812 8084
rect 314752 8032 314804 8084
rect 405372 8032 405424 8084
rect 552664 8032 552716 8084
rect 30104 7896 30156 7948
rect 243084 7896 243136 7948
rect 251180 7896 251232 7948
rect 314844 7964 314896 8016
rect 406752 7964 406804 8016
rect 556160 7964 556212 8016
rect 26516 7828 26568 7880
rect 242992 7828 243044 7880
rect 254676 7828 254728 7880
rect 313372 7896 313424 7948
rect 408224 7896 408276 7948
rect 559748 7896 559800 7948
rect 312084 7828 312136 7880
rect 409512 7828 409564 7880
rect 563244 7828 563296 7880
rect 21824 7760 21876 7812
rect 241796 7760 241848 7812
rect 247592 7760 247644 7812
rect 310612 7760 310664 7812
rect 410984 7760 411036 7812
rect 566832 7760 566884 7812
rect 17040 7692 17092 7744
rect 240140 7692 240192 7744
rect 244096 7692 244148 7744
rect 309324 7692 309376 7744
rect 410892 7692 410944 7744
rect 570328 7692 570380 7744
rect 12348 7624 12400 7676
rect 237380 7624 237432 7676
rect 240508 7624 240560 7676
rect 309232 7624 309284 7676
rect 412272 7624 412324 7676
rect 573916 7624 573968 7676
rect 4068 7556 4120 7608
rect 236184 7556 236236 7608
rect 237012 7556 237064 7608
rect 307852 7556 307904 7608
rect 413744 7556 413796 7608
rect 577412 7556 577464 7608
rect 141240 7488 141292 7540
rect 277492 7488 277544 7540
rect 371056 7488 371108 7540
rect 144736 7420 144788 7472
rect 278964 7420 279016 7472
rect 369676 7420 369728 7472
rect 148324 7352 148376 7404
rect 280344 7352 280396 7404
rect 368204 7352 368256 7404
rect 432052 7352 432104 7404
rect 151820 7284 151872 7336
rect 281724 7284 281776 7336
rect 368296 7284 368348 7336
rect 155408 7216 155460 7268
rect 283012 7216 283064 7268
rect 367008 7216 367060 7268
rect 424968 7216 425020 7268
rect 425704 7284 425756 7336
rect 427268 7284 427320 7336
rect 435364 7488 435416 7540
rect 437940 7488 437992 7540
rect 439136 7352 439188 7404
rect 435548 7284 435600 7336
rect 428464 7216 428516 7268
rect 158904 7148 158956 7200
rect 283104 7148 283156 7200
rect 365536 7148 365588 7200
rect 421380 7148 421432 7200
rect 229836 7080 229888 7132
rect 305092 7080 305144 7132
rect 364156 7080 364208 7132
rect 417884 7080 417936 7132
rect 233424 7012 233476 7064
rect 306564 7012 306616 7064
rect 362592 7012 362644 7064
rect 414296 7012 414348 7064
rect 234620 6808 234672 6860
rect 580172 6808 580224 6860
rect 169576 6740 169628 6792
rect 287244 6740 287296 6792
rect 382096 6740 382148 6792
rect 476948 6740 477000 6792
rect 166080 6672 166132 6724
rect 285864 6672 285916 6724
rect 384856 6672 384908 6724
rect 481732 6672 481784 6724
rect 130568 6604 130620 6656
rect 274824 6604 274876 6656
rect 384764 6604 384816 6656
rect 485228 6604 485280 6656
rect 69112 6536 69164 6588
rect 255412 6536 255464 6588
rect 386328 6536 386380 6588
rect 488816 6536 488868 6588
rect 65524 6468 65576 6520
rect 254032 6468 254084 6520
rect 387708 6468 387760 6520
rect 492312 6468 492364 6520
rect 62028 6400 62080 6452
rect 254124 6400 254176 6452
rect 389088 6400 389140 6452
rect 495900 6400 495952 6452
rect 58440 6332 58492 6384
rect 252652 6332 252704 6384
rect 299664 6332 299716 6384
rect 316684 6332 316736 6384
rect 390192 6332 390244 6384
rect 499396 6332 499448 6384
rect 54944 6264 54996 6316
rect 251364 6264 251416 6316
rect 259460 6264 259512 6316
rect 295984 6264 296036 6316
rect 303160 6264 303212 6316
rect 327724 6264 327776 6316
rect 390376 6264 390428 6316
rect 502892 6264 502944 6316
rect 51356 6196 51408 6248
rect 250076 6196 250128 6248
rect 268844 6196 268896 6248
rect 317696 6196 317748 6248
rect 371884 6196 371936 6248
rect 378876 6196 378928 6248
rect 391664 6196 391716 6248
rect 506572 6196 506624 6248
rect 47860 6128 47912 6180
rect 248512 6128 248564 6180
rect 257068 6128 257120 6180
rect 313280 6128 313332 6180
rect 370504 6128 370556 6180
rect 385960 6128 386012 6180
rect 393136 6128 393188 6180
rect 510068 6128 510120 6180
rect 173164 6060 173216 6112
rect 287152 6060 287204 6112
rect 382004 6060 382056 6112
rect 473452 6060 473504 6112
rect 176660 5992 176712 6044
rect 288624 5992 288676 6044
rect 380716 5992 380768 6044
rect 469864 5992 469916 6044
rect 180248 5924 180300 5976
rect 290004 5924 290056 5976
rect 379428 5924 379480 5976
rect 466276 5924 466328 5976
rect 468484 5924 468536 5976
rect 474556 5924 474608 5976
rect 183744 5856 183796 5908
rect 291384 5856 291436 5908
rect 377956 5856 378008 5908
rect 462780 5856 462832 5908
rect 187332 5788 187384 5840
rect 292672 5788 292724 5840
rect 377864 5788 377916 5840
rect 459192 5788 459244 5840
rect 190828 5720 190880 5772
rect 292764 5720 292816 5772
rect 376668 5720 376720 5772
rect 455696 5720 455748 5772
rect 194416 5652 194468 5704
rect 294236 5652 294288 5704
rect 375196 5652 375248 5704
rect 452108 5652 452160 5704
rect 363604 5516 363656 5568
rect 367008 5516 367060 5568
rect 475384 5516 475436 5568
rect 480536 5516 480588 5568
rect 486516 5516 486568 5568
rect 487620 5516 487672 5568
rect 497464 5516 497516 5568
rect 498200 5516 498252 5568
rect 504364 5516 504416 5568
rect 505376 5516 505428 5568
rect 186228 5448 186280 5500
rect 215944 5448 215996 5500
rect 218060 5448 218112 5500
rect 302332 5448 302384 5500
rect 355784 5448 355836 5500
rect 391848 5448 391900 5500
rect 402704 5448 402756 5500
rect 540796 5448 540848 5500
rect 189724 5380 189776 5432
rect 214288 5380 214340 5432
rect 214472 5380 214524 5432
rect 301044 5380 301096 5432
rect 357256 5380 357308 5432
rect 395344 5380 395396 5432
rect 404176 5380 404228 5432
rect 544384 5380 544436 5432
rect 210976 5312 211028 5364
rect 299756 5312 299808 5364
rect 358544 5312 358596 5364
rect 400128 5312 400180 5364
rect 404084 5312 404136 5364
rect 547880 5312 547932 5364
rect 136456 5244 136508 5296
rect 204904 5244 204956 5296
rect 207388 5244 207440 5296
rect 298284 5244 298336 5296
rect 358636 5244 358688 5296
rect 398932 5244 398984 5296
rect 405556 5244 405608 5296
rect 551468 5244 551520 5296
rect 203892 5176 203944 5228
rect 296904 5176 296956 5228
rect 359832 5176 359884 5228
rect 402520 5176 402572 5228
rect 406844 5176 406896 5228
rect 554964 5176 555016 5228
rect 132960 5108 133012 5160
rect 274640 5108 274692 5160
rect 278320 5108 278372 5160
rect 320364 5108 320416 5160
rect 359924 5108 359976 5160
rect 403624 5108 403676 5160
rect 408316 5108 408368 5160
rect 558552 5108 558604 5160
rect 129372 5040 129424 5092
rect 274732 5040 274784 5092
rect 274824 5040 274876 5092
rect 318892 5040 318944 5092
rect 361212 5040 361264 5092
rect 406016 5040 406068 5092
rect 409604 5040 409656 5092
rect 409696 5040 409748 5092
rect 562048 5040 562100 5092
rect 7656 4972 7708 5024
rect 236092 4972 236144 5024
rect 246396 4972 246448 5024
rect 310520 4972 310572 5024
rect 361304 4972 361356 5024
rect 407212 4972 407264 5024
rect 565636 4972 565688 5024
rect 2872 4904 2924 4956
rect 234804 4904 234856 4956
rect 242900 4904 242952 4956
rect 309140 4904 309192 4956
rect 361396 4904 361448 4956
rect 409604 4904 409656 4956
rect 411076 4904 411128 4956
rect 569132 4904 569184 4956
rect 1676 4836 1728 4888
rect 234896 4836 234948 4888
rect 239312 4836 239364 4888
rect 307760 4836 307812 4888
rect 362684 4836 362736 4888
rect 410800 4836 410852 4888
rect 412364 4836 412416 4888
rect 572720 4836 572772 4888
rect 572 4768 624 4820
rect 234712 4768 234764 4820
rect 235816 4768 235868 4820
rect 306472 4768 306524 4820
rect 362776 4768 362828 4820
rect 413100 4768 413152 4820
rect 413836 4768 413888 4820
rect 576308 4768 576360 4820
rect 193220 4700 193272 4752
rect 220084 4700 220136 4752
rect 221556 4700 221608 4752
rect 302516 4700 302568 4752
rect 355876 4700 355928 4752
rect 388260 4700 388312 4752
rect 401324 4700 401376 4752
rect 537208 4700 537260 4752
rect 171968 4632 172020 4684
rect 222844 4632 222896 4684
rect 225144 4632 225196 4684
rect 303804 4632 303856 4684
rect 354496 4632 354548 4684
rect 384764 4632 384816 4684
rect 399852 4632 399904 4684
rect 533712 4632 533764 4684
rect 228732 4564 228784 4616
rect 305000 4564 305052 4616
rect 353116 4564 353168 4616
rect 381176 4564 381228 4616
rect 398656 4564 398708 4616
rect 530124 4564 530176 4616
rect 232228 4496 232280 4548
rect 306380 4496 306432 4548
rect 351736 4496 351788 4548
rect 377680 4496 377732 4548
rect 398564 4496 398616 4548
rect 526628 4496 526680 4548
rect 281908 4428 281960 4480
rect 321744 4428 321796 4480
rect 350264 4428 350316 4480
rect 374092 4428 374144 4480
rect 397092 4428 397144 4480
rect 523040 4428 523092 4480
rect 285404 4360 285456 4412
rect 323032 4360 323084 4412
rect 395804 4360 395856 4412
rect 519544 4360 519596 4412
rect 288992 4292 289044 4344
rect 323124 4292 323176 4344
rect 394424 4292 394476 4344
rect 515956 4292 516008 4344
rect 200304 4224 200356 4276
rect 208952 4224 209004 4276
rect 292580 4224 292632 4276
rect 324596 4224 324648 4276
rect 332600 4224 332652 4276
rect 332784 4224 332836 4276
rect 392952 4224 393004 4276
rect 512460 4224 512512 4276
rect 143540 4156 143592 4208
rect 144828 4156 144880 4208
rect 184940 4156 184992 4208
rect 186136 4156 186188 4208
rect 201500 4156 201552 4208
rect 202788 4156 202840 4208
rect 226340 4156 226392 4208
rect 227628 4156 227680 4208
rect 388444 4156 388496 4208
rect 393044 4156 393096 4208
rect 418804 4156 418856 4208
rect 420184 4156 420236 4208
rect 11152 4088 11204 4140
rect 18604 4088 18656 4140
rect 34796 4088 34848 4140
rect 36544 4088 36596 4140
rect 82084 4020 82136 4072
rect 259736 4088 259788 4140
rect 306748 4088 306800 4140
rect 328552 4088 328604 4140
rect 343548 4088 343600 4140
rect 350448 4088 350500 4140
rect 351828 4088 351880 4140
rect 375288 4088 375340 4140
rect 402796 4088 402848 4140
rect 258172 4020 258224 4072
rect 309048 4020 309100 4072
rect 330116 4020 330168 4072
rect 332692 4020 332744 4072
rect 336004 4020 336056 4072
rect 343456 4020 343508 4072
rect 348056 4020 348108 4072
rect 350356 4020 350408 4072
rect 372896 4020 372948 4072
rect 402612 4020 402664 4072
rect 543188 4020 543240 4072
rect 43076 3952 43128 4004
rect 51724 3952 51776 4004
rect 53656 3952 53708 4004
rect 57244 3952 57296 4004
rect 75000 3952 75052 4004
rect 258080 3952 258132 4004
rect 305552 3952 305604 4004
rect 328736 3952 328788 4004
rect 329196 3952 329248 4004
rect 335544 3952 335596 4004
rect 342168 3952 342220 4004
rect 346952 3952 347004 4004
rect 353208 3952 353260 4004
rect 379980 3952 380032 4004
rect 404268 3952 404320 4004
rect 546684 3952 546736 4004
rect 38384 3884 38436 3936
rect 47584 3884 47636 3936
rect 50160 3884 50212 3936
rect 68284 3884 68336 3936
rect 71504 3884 71556 3936
rect 256700 3884 256752 3936
rect 301964 3884 302016 3936
rect 5264 3816 5316 3868
rect 7564 3816 7616 3868
rect 41880 3816 41932 3868
rect 54484 3816 54536 3868
rect 67916 3816 67968 3868
rect 255320 3816 255372 3868
rect 297272 3816 297324 3868
rect 325792 3884 325844 3936
rect 326804 3884 326856 3936
rect 335636 3884 335688 3936
rect 344284 3884 344336 3936
rect 351644 3884 351696 3936
rect 354588 3884 354640 3936
rect 387156 3884 387208 3936
rect 405648 3884 405700 3936
rect 550272 3884 550324 3936
rect 320916 3816 320968 3868
rect 329104 3816 329156 3868
rect 333888 3816 333940 3868
rect 336924 3816 336976 3868
rect 345756 3816 345808 3868
rect 356336 3816 356388 3868
rect 357348 3816 357400 3868
rect 35992 3748 36044 3800
rect 50344 3748 50396 3800
rect 64328 3748 64380 3800
rect 253940 3748 253992 3800
rect 293684 3748 293736 3800
rect 327264 3748 327316 3800
rect 334072 3748 334124 3800
rect 343364 3748 343416 3800
rect 349252 3748 349304 3800
rect 355968 3748 356020 3800
rect 358728 3748 358780 3800
rect 390652 3816 390704 3868
rect 406936 3816 406988 3868
rect 553768 3816 553820 3868
rect 394240 3748 394292 3800
rect 407028 3748 407080 3800
rect 557356 3748 557408 3800
rect 23020 3680 23072 3732
rect 39304 3680 39356 3732
rect 20628 3612 20680 3664
rect 43444 3680 43496 3732
rect 45376 3680 45428 3732
rect 58624 3680 58676 3732
rect 60832 3680 60884 3732
rect 252836 3680 252888 3732
rect 291384 3680 291436 3732
rect 324320 3680 324372 3732
rect 324412 3680 324464 3732
rect 334164 3680 334216 3732
rect 346308 3680 346360 3732
rect 39580 3612 39632 3664
rect 18236 3544 18288 3596
rect 28908 3544 28960 3596
rect 35164 3544 35216 3596
rect 40684 3544 40736 3596
rect 41328 3544 41380 3596
rect 48964 3544 49016 3596
rect 49608 3544 49660 3596
rect 52552 3544 52604 3596
rect 53748 3544 53800 3596
rect 248696 3612 248748 3664
rect 284300 3612 284352 3664
rect 321836 3612 321888 3664
rect 247224 3544 247276 3596
rect 279516 3544 279568 3596
rect 32312 3476 32364 3528
rect 32404 3476 32456 3528
rect 244464 3476 244516 3528
rect 249984 3476 250036 3528
rect 251088 3476 251140 3528
rect 255872 3476 255924 3528
rect 256608 3476 256660 3528
rect 262956 3476 263008 3528
rect 263508 3476 263560 3528
rect 264152 3476 264204 3528
rect 264888 3476 264940 3528
rect 266544 3476 266596 3528
rect 267648 3476 267700 3528
rect 271236 3476 271288 3528
rect 271788 3476 271840 3528
rect 273628 3476 273680 3528
rect 274548 3476 274600 3528
rect 276020 3476 276072 3528
rect 277308 3476 277360 3528
rect 280712 3476 280764 3528
rect 281448 3476 281500 3528
rect 286600 3544 286652 3596
rect 324504 3612 324556 3664
rect 325608 3612 325660 3664
rect 335452 3612 335504 3664
rect 347136 3612 347188 3664
rect 397736 3680 397788 3732
rect 408408 3680 408460 3732
rect 560852 3680 560904 3732
rect 320272 3476 320324 3528
rect 323216 3544 323268 3596
rect 323308 3544 323360 3596
rect 332600 3544 332652 3596
rect 342076 3544 342128 3596
rect 344560 3544 344612 3596
rect 347596 3544 347648 3596
rect 358728 3612 358780 3664
rect 360016 3612 360068 3664
rect 401324 3612 401376 3664
rect 409788 3612 409840 3664
rect 564440 3612 564492 3664
rect 322112 3476 322164 3528
rect 13544 3408 13596 3460
rect 22744 3408 22796 3460
rect 25320 3408 25372 3460
rect 241612 3408 241664 3460
rect 267740 3408 267792 3460
rect 269028 3408 269080 3460
rect 272432 3408 272484 3460
rect 318984 3408 319036 3460
rect 319720 3408 319772 3460
rect 19432 3340 19484 3392
rect 25504 3340 25556 3392
rect 31300 3340 31352 3392
rect 33784 3340 33836 3392
rect 44272 3340 44324 3392
rect 45468 3340 45520 3392
rect 46664 3340 46716 3392
rect 56048 3340 56100 3392
rect 56508 3340 56560 3392
rect 59636 3340 59688 3392
rect 60648 3340 60700 3392
rect 66720 3340 66772 3392
rect 67548 3340 67600 3392
rect 73804 3340 73856 3392
rect 74448 3340 74500 3392
rect 77392 3340 77444 3392
rect 78588 3340 78640 3392
rect 80888 3340 80940 3392
rect 81348 3340 81400 3392
rect 78588 3204 78640 3256
rect 84476 3340 84528 3392
rect 87604 3340 87656 3392
rect 90364 3340 90416 3392
rect 91008 3340 91060 3392
rect 91560 3340 91612 3392
rect 93124 3340 93176 3392
rect 83280 3272 83332 3324
rect 84108 3272 84160 3324
rect 87972 3272 88024 3324
rect 88984 3272 89036 3324
rect 261024 3340 261076 3392
rect 287796 3340 287848 3392
rect 288348 3340 288400 3392
rect 296076 3340 296128 3392
rect 296628 3340 296680 3392
rect 298468 3340 298520 3392
rect 299388 3340 299440 3392
rect 307944 3340 307996 3392
rect 329840 3340 329892 3392
rect 331588 3476 331640 3528
rect 332508 3476 332560 3528
rect 337476 3476 337528 3528
rect 338120 3476 338172 3528
rect 345664 3476 345716 3528
rect 352840 3476 352892 3528
rect 359924 3544 359976 3596
rect 360108 3544 360160 3596
rect 404820 3544 404872 3596
rect 411168 3544 411220 3596
rect 568028 3544 568080 3596
rect 361120 3476 361172 3528
rect 361488 3476 361540 3528
rect 408408 3476 408460 3528
rect 412548 3476 412600 3528
rect 571524 3476 571576 3528
rect 330392 3408 330444 3460
rect 333244 3408 333296 3460
rect 335084 3408 335136 3460
rect 338212 3408 338264 3460
rect 347688 3408 347740 3460
rect 362316 3408 362368 3460
rect 362868 3408 362920 3460
rect 411904 3408 411956 3460
rect 412456 3408 412508 3460
rect 575112 3408 575164 3460
rect 334348 3340 334400 3392
rect 350540 3340 350592 3392
rect 371700 3340 371752 3392
rect 382188 3340 382240 3392
rect 475752 3340 475804 3392
rect 481640 3340 481692 3392
rect 482836 3340 482888 3392
rect 489184 3340 489236 3392
rect 489920 3340 489972 3392
rect 85672 3204 85724 3256
rect 93952 3272 94004 3324
rect 95056 3272 95108 3324
rect 97448 3272 97500 3324
rect 97908 3272 97960 3324
rect 98644 3272 98696 3324
rect 99288 3272 99340 3324
rect 101036 3272 101088 3324
rect 102048 3272 102100 3324
rect 262496 3272 262548 3324
rect 310244 3272 310296 3324
rect 330024 3272 330076 3324
rect 348976 3272 349028 3324
rect 369400 3272 369452 3324
rect 380808 3272 380860 3324
rect 468668 3272 468720 3324
rect 485044 3272 485096 3324
rect 502984 3272 503036 3324
rect 504180 3272 504232 3324
rect 506480 3272 506532 3324
rect 507676 3272 507728 3324
rect 515404 3272 515456 3324
rect 517152 3272 517204 3324
rect 519636 3272 519688 3324
rect 521844 3272 521896 3324
rect 522304 3272 522356 3324
rect 524236 3272 524288 3324
rect 530584 3340 530636 3392
rect 531320 3340 531372 3392
rect 533344 3340 533396 3392
rect 534908 3340 534960 3392
rect 539600 3340 539652 3392
rect 540244 3340 540296 3392
rect 541992 3340 542044 3392
rect 532516 3272 532568 3324
rect 92756 3204 92808 3256
rect 262312 3204 262364 3256
rect 312636 3204 312688 3256
rect 331404 3204 331456 3256
rect 349068 3204 349120 3256
rect 365812 3204 365864 3256
rect 377772 3204 377824 3256
rect 461584 3204 461636 3256
rect 526444 3204 526496 3256
rect 527824 3204 527876 3256
rect 57244 3136 57296 3188
rect 61384 3136 61436 3188
rect 89168 3136 89220 3188
rect 96252 3068 96304 3120
rect 263784 3136 263836 3188
rect 311440 3136 311492 3188
rect 329932 3136 329984 3188
rect 349804 3136 349856 3188
rect 102232 3068 102284 3120
rect 104164 3068 104216 3120
rect 105728 3068 105780 3120
rect 106188 3068 106240 3120
rect 106924 3068 106976 3120
rect 107568 3068 107620 3120
rect 108120 3068 108172 3120
rect 108948 3068 109000 3120
rect 109316 3068 109368 3120
rect 111064 3068 111116 3120
rect 265256 3068 265308 3120
rect 313832 3068 313884 3120
rect 331496 3068 331548 3120
rect 338672 3068 338724 3120
rect 339592 3068 339644 3120
rect 347044 3068 347096 3120
rect 354036 3068 354088 3120
rect 355232 3136 355284 3188
rect 357532 3068 357584 3120
rect 358084 3068 358136 3120
rect 363512 3068 363564 3120
rect 27712 3000 27764 3052
rect 29644 3000 29696 3052
rect 103336 3000 103388 3052
rect 266636 3000 266688 3052
rect 317328 3000 317380 3052
rect 332968 3000 333020 3052
rect 348424 3000 348476 3052
rect 99840 2932 99892 2984
rect 9956 2864 10008 2916
rect 14464 2864 14516 2916
rect 110512 2932 110564 2984
rect 267924 2932 267976 2984
rect 304356 2932 304408 2984
rect 304908 2932 304960 2984
rect 315028 2932 315080 2984
rect 331680 2932 331732 2984
rect 336280 2932 336332 2984
rect 338304 2932 338356 2984
rect 348516 2932 348568 2984
rect 364616 3136 364668 3188
rect 375196 3136 375248 3188
rect 454500 3136 454552 3188
rect 512644 3136 512696 3188
rect 513564 3136 513616 3188
rect 373908 3068 373960 3120
rect 447416 3068 447468 3120
rect 371148 3000 371200 3052
rect 440240 3000 440292 3052
rect 440332 3000 440384 3052
rect 441528 3000 441580 3052
rect 369768 2932 369820 2984
rect 433248 2932 433300 2984
rect 114008 2864 114060 2916
rect 114468 2864 114520 2916
rect 115204 2864 115256 2916
rect 115848 2864 115900 2916
rect 116400 2864 116452 2916
rect 117228 2864 117280 2916
rect 118792 2864 118844 2916
rect 119804 2864 119856 2916
rect 117596 2796 117648 2848
rect 122288 2864 122340 2916
rect 122748 2864 122800 2916
rect 123484 2864 123536 2916
rect 124128 2864 124180 2916
rect 124680 2864 124732 2916
rect 125416 2864 125468 2916
rect 121092 2796 121144 2848
rect 270776 2864 270828 2916
rect 316224 2864 316276 2916
rect 331312 2864 331364 2916
rect 365628 2864 365680 2916
rect 422576 2864 422628 2916
rect 272064 2796 272116 2848
rect 318524 2796 318576 2848
rect 332784 2796 332836 2848
rect 364248 2796 364300 2848
rect 415492 2796 415544 2848
rect 168380 1640 168432 1692
rect 169668 1640 169720 1692
rect 456800 1368 456852 1420
rect 458088 1368 458140 1420
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 89364 703582 89668 703610
rect 8128 700330 8156 703520
rect 8116 700324 8168 700330
rect 8116 700266 8168 700272
rect 24320 699718 24348 703520
rect 40512 700466 40540 703520
rect 40500 700460 40552 700466
rect 40500 700402 40552 700408
rect 41328 700460 41380 700466
rect 41328 700402 41380 700408
rect 24308 699712 24360 699718
rect 24308 699654 24360 699660
rect 24768 699712 24820 699718
rect 24768 699654 24820 699660
rect 3422 684312 3478 684321
rect 3422 684247 3478 684256
rect 3330 619168 3386 619177
rect 3330 619103 3386 619112
rect 3344 618322 3372 619103
rect 3332 618316 3384 618322
rect 3332 618258 3384 618264
rect 3330 606112 3386 606121
rect 3330 606047 3386 606056
rect 3344 605878 3372 606047
rect 3332 605872 3384 605878
rect 3332 605814 3384 605820
rect 3054 566944 3110 566953
rect 3054 566879 3110 566888
rect 3068 565894 3096 566879
rect 3056 565888 3108 565894
rect 3056 565830 3108 565836
rect 3330 553888 3386 553897
rect 3330 553823 3386 553832
rect 3344 553450 3372 553823
rect 3332 553444 3384 553450
rect 3332 553386 3384 553392
rect 3330 514856 3386 514865
rect 3330 514791 3332 514800
rect 3384 514791 3386 514800
rect 3332 514762 3384 514768
rect 3238 501800 3294 501809
rect 3238 501735 3294 501744
rect 3252 501022 3280 501735
rect 3240 501016 3292 501022
rect 3240 500958 3292 500964
rect 3436 460494 3464 684247
rect 3514 671256 3570 671265
rect 3514 671191 3570 671200
rect 3528 670750 3556 671191
rect 3516 670744 3568 670750
rect 3516 670686 3568 670692
rect 3514 658200 3570 658209
rect 3514 658135 3570 658144
rect 3528 656946 3556 658135
rect 3516 656940 3568 656946
rect 3516 656882 3568 656888
rect 3514 632088 3570 632097
rect 3514 632023 3570 632032
rect 3528 465746 3556 632023
rect 3606 580000 3662 580009
rect 3606 579935 3662 579944
rect 3620 465882 3648 579935
rect 3698 527912 3754 527921
rect 3698 527847 3754 527856
rect 3712 466018 3740 527847
rect 3882 475688 3938 475697
rect 3882 475623 3938 475632
rect 3712 465990 3832 466018
rect 3620 465854 3740 465882
rect 3528 465718 3648 465746
rect 3514 462632 3570 462641
rect 3514 462567 3570 462576
rect 3528 462398 3556 462567
rect 3516 462392 3568 462398
rect 3516 462334 3568 462340
rect 3424 460488 3476 460494
rect 3424 460430 3476 460436
rect 3620 460426 3648 465718
rect 3608 460420 3660 460426
rect 3608 460362 3660 460368
rect 3712 460358 3740 465854
rect 3700 460352 3752 460358
rect 3700 460294 3752 460300
rect 3804 460290 3832 465990
rect 3792 460284 3844 460290
rect 3792 460226 3844 460232
rect 3896 460222 3924 475623
rect 24780 460562 24808 699654
rect 41340 460630 41368 700402
rect 72988 700398 73016 703520
rect 89180 703474 89208 703520
rect 89364 703474 89392 703582
rect 89180 703446 89392 703474
rect 72976 700392 73028 700398
rect 72976 700334 73028 700340
rect 89640 460698 89668 703582
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 154316 703582 154528 703610
rect 105464 700534 105492 703520
rect 137848 700670 137876 703520
rect 154132 703474 154160 703520
rect 154316 703474 154344 703582
rect 154132 703446 154344 703474
rect 137836 700664 137888 700670
rect 137836 700606 137888 700612
rect 105452 700528 105504 700534
rect 105452 700470 105504 700476
rect 106188 700528 106240 700534
rect 106188 700470 106240 700476
rect 106200 460766 106228 700470
rect 154500 460834 154528 703582
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 284036 703582 284248 703610
rect 170324 699718 170352 703520
rect 202800 700942 202828 703520
rect 218992 702434 219020 703520
rect 218992 702406 219388 702434
rect 202788 700936 202840 700942
rect 202788 700878 202840 700884
rect 170312 699712 170364 699718
rect 170312 699654 170364 699660
rect 171048 699712 171100 699718
rect 171048 699654 171100 699660
rect 171060 460902 171088 699654
rect 171048 460896 171100 460902
rect 171048 460838 171100 460844
rect 154488 460828 154540 460834
rect 154488 460770 154540 460776
rect 106188 460760 106240 460766
rect 106188 460702 106240 460708
rect 89628 460692 89680 460698
rect 89628 460634 89680 460640
rect 41328 460624 41380 460630
rect 41328 460566 41380 460572
rect 24768 460556 24820 460562
rect 24768 460498 24820 460504
rect 3884 460216 3936 460222
rect 3884 460158 3936 460164
rect 219360 460154 219388 702406
rect 235184 699718 235212 703520
rect 267660 700126 267688 703520
rect 283852 703474 283880 703520
rect 284036 703474 284064 703582
rect 283852 703446 284064 703474
rect 267648 700120 267700 700126
rect 267648 700062 267700 700068
rect 235172 699712 235224 699718
rect 235172 699654 235224 699660
rect 235908 699712 235960 699718
rect 235908 699654 235960 699660
rect 219348 460148 219400 460154
rect 219348 460090 219400 460096
rect 235920 460086 235948 699654
rect 235908 460080 235960 460086
rect 235908 460022 235960 460028
rect 284220 460018 284248 703582
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 300136 699718 300164 703520
rect 317328 701004 317380 701010
rect 317328 700946 317380 700952
rect 313188 700868 313240 700874
rect 313188 700810 313240 700816
rect 311808 700732 311860 700738
rect 311808 700674 311860 700680
rect 309048 700596 309100 700602
rect 309048 700538 309100 700544
rect 307668 700460 307720 700466
rect 307668 700402 307720 700408
rect 300124 699712 300176 699718
rect 300124 699654 300176 699660
rect 300768 699712 300820 699718
rect 300768 699654 300820 699660
rect 299388 643136 299440 643142
rect 299388 643078 299440 643084
rect 298008 616888 298060 616894
rect 298008 616830 298060 616836
rect 295248 590708 295300 590714
rect 295248 590650 295300 590656
rect 293868 563100 293920 563106
rect 293868 563042 293920 563048
rect 289728 536852 289780 536858
rect 289728 536794 289780 536800
rect 288348 510672 288400 510678
rect 288348 510614 288400 510620
rect 285588 484424 285640 484430
rect 285588 484366 285640 484372
rect 284208 460012 284260 460018
rect 284208 459954 284260 459960
rect 281448 459808 281500 459814
rect 281448 459750 281500 459756
rect 272340 459672 272392 459678
rect 272340 459614 272392 459620
rect 267464 459604 267516 459610
rect 267464 459546 267516 459552
rect 231124 458788 231176 458794
rect 231124 458730 231176 458736
rect 222844 458652 222896 458658
rect 222844 458594 222896 458600
rect 3424 458244 3476 458250
rect 3424 458186 3476 458192
rect 3332 449880 3384 449886
rect 3332 449822 3384 449828
rect 3344 449585 3372 449822
rect 3330 449576 3386 449585
rect 3330 449511 3386 449520
rect 3436 423609 3464 458186
rect 4804 456816 4856 456822
rect 4804 456758 4856 456764
rect 3422 423600 3478 423609
rect 3422 423535 3478 423544
rect 3424 411256 3476 411262
rect 3424 411198 3476 411204
rect 3436 410553 3464 411198
rect 3422 410544 3478 410553
rect 3422 410479 3478 410488
rect 3240 398812 3292 398818
rect 3240 398754 3292 398760
rect 3252 397497 3280 398754
rect 3238 397488 3294 397497
rect 3238 397423 3294 397432
rect 4816 371482 4844 456758
rect 222856 411262 222884 458594
rect 228364 458380 228416 458386
rect 228364 458322 228416 458328
rect 226984 457224 227036 457230
rect 226984 457166 227036 457172
rect 224224 457088 224276 457094
rect 224224 457030 224276 457036
rect 222844 411256 222896 411262
rect 222844 411198 222896 411204
rect 2780 371476 2832 371482
rect 2780 371418 2832 371424
rect 4804 371476 4856 371482
rect 4804 371418 4856 371424
rect 2792 371385 2820 371418
rect 2778 371376 2834 371385
rect 2778 371311 2834 371320
rect 224236 358766 224264 457030
rect 3332 358760 3384 358766
rect 3332 358702 3384 358708
rect 224224 358760 224276 358766
rect 224224 358702 224276 358708
rect 3344 358465 3372 358702
rect 3330 358456 3386 358465
rect 3330 358391 3386 358400
rect 226996 346390 227024 457166
rect 3148 346384 3200 346390
rect 3148 346326 3200 346332
rect 226984 346384 227036 346390
rect 226984 346326 227036 346332
rect 3160 345409 3188 346326
rect 3146 345400 3202 345409
rect 3146 345335 3202 345344
rect 220084 336728 220136 336734
rect 220084 336670 220136 336676
rect 215944 336660 215996 336666
rect 215944 336602 215996 336608
rect 214564 336592 214616 336598
rect 214564 336534 214616 336540
rect 209044 336524 209096 336530
rect 209044 336466 209096 336472
rect 125508 336456 125560 336462
rect 43442 336424 43498 336433
rect 125508 336398 125560 336404
rect 43442 336359 43498 336368
rect 114468 336388 114520 336394
rect 25502 336288 25558 336297
rect 25502 336223 25558 336232
rect 18602 336152 18658 336161
rect 18602 336087 18658 336096
rect 7562 336016 7618 336025
rect 7562 335951 7618 335960
rect 3422 320104 3478 320113
rect 3422 320039 3478 320048
rect 3436 319297 3464 320039
rect 3422 319288 3478 319297
rect 3422 319223 3478 319232
rect 3330 293856 3386 293865
rect 3330 293791 3386 293800
rect 3344 293185 3372 293791
rect 3330 293176 3386 293185
rect 3330 293111 3386 293120
rect 3422 255232 3478 255241
rect 3422 255167 3478 255176
rect 3436 254153 3464 255167
rect 3422 254144 3478 254153
rect 3422 254079 3478 254088
rect 3332 215280 3384 215286
rect 3332 215222 3384 215228
rect 3344 214985 3372 215222
rect 3330 214976 3386 214985
rect 3330 214911 3386 214920
rect 3422 202872 3478 202881
rect 3422 202807 3478 202816
rect 3436 201929 3464 202807
rect 3422 201920 3478 201929
rect 3422 201855 3478 201864
rect 3422 164112 3478 164121
rect 3422 164047 3478 164056
rect 3436 162897 3464 164047
rect 3422 162888 3478 162897
rect 3422 162823 3478 162832
rect 3422 138000 3478 138009
rect 3422 137935 3478 137944
rect 3436 136785 3464 137935
rect 3422 136776 3478 136785
rect 3422 136711 3478 136720
rect 3422 111752 3478 111761
rect 3422 111687 3478 111696
rect 3436 110673 3464 111687
rect 3422 110664 3478 110673
rect 3422 110599 3478 110608
rect 3422 85504 3478 85513
rect 3422 85439 3478 85448
rect 3436 84697 3464 85439
rect 3422 84688 3478 84697
rect 3422 84623 3478 84632
rect 3330 59256 3386 59265
rect 3330 59191 3386 59200
rect 3344 58585 3372 59191
rect 3330 58576 3386 58585
rect 3330 58511 3386 58520
rect 3424 45552 3476 45558
rect 3422 45520 3424 45529
rect 3476 45520 3478 45529
rect 3422 45455 3478 45464
rect 3330 33144 3386 33153
rect 3330 33079 3386 33088
rect 3344 32473 3372 33079
rect 3330 32464 3386 32473
rect 3330 32399 3386 32408
rect 3424 20664 3476 20670
rect 3424 20606 3476 20612
rect 3436 19417 3464 20606
rect 3422 19408 3478 19417
rect 3422 19343 3478 19352
rect 4068 7608 4120 7614
rect 4068 7550 4120 7556
rect 2872 4956 2924 4962
rect 2872 4898 2924 4904
rect 1676 4888 1728 4894
rect 1676 4830 1728 4836
rect 572 4820 624 4826
rect 572 4762 624 4768
rect 584 480 612 4762
rect 1688 480 1716 4830
rect 2884 480 2912 4898
rect 4080 480 4108 7550
rect 7576 3874 7604 335951
rect 14464 327752 14516 327758
rect 14464 327694 14516 327700
rect 8760 8968 8812 8974
rect 8760 8910 8812 8916
rect 7656 5024 7708 5030
rect 7656 4966 7708 4972
rect 5264 3868 5316 3874
rect 5264 3810 5316 3816
rect 7564 3868 7616 3874
rect 7564 3810 7616 3816
rect 5276 480 5304 3810
rect 6458 3360 6514 3369
rect 6458 3295 6514 3304
rect 6472 480 6500 3295
rect 7668 480 7696 4966
rect 8772 480 8800 8910
rect 12348 7676 12400 7682
rect 12348 7618 12400 7624
rect 11152 4140 11204 4146
rect 11152 4082 11204 4088
rect 9956 2916 10008 2922
rect 9956 2858 10008 2864
rect 9968 480 9996 2858
rect 11164 480 11192 4082
rect 12360 480 12388 7618
rect 13544 3460 13596 3466
rect 13544 3402 13596 3408
rect 13556 480 13584 3402
rect 14476 2922 14504 327694
rect 17040 7744 17092 7750
rect 17040 7686 17092 7692
rect 15934 3632 15990 3641
rect 15934 3567 15990 3576
rect 14738 3496 14794 3505
rect 14738 3431 14794 3440
rect 14464 2916 14516 2922
rect 14464 2858 14516 2864
rect 14752 480 14780 3431
rect 15948 480 15976 3567
rect 17052 480 17080 7686
rect 18616 4146 18644 336087
rect 22744 334620 22796 334626
rect 22744 334562 22796 334568
rect 21824 7812 21876 7818
rect 21824 7754 21876 7760
rect 18604 4140 18656 4146
rect 18604 4082 18656 4088
rect 20628 3664 20680 3670
rect 20628 3606 20680 3612
rect 18236 3596 18288 3602
rect 18236 3538 18288 3544
rect 18248 480 18276 3538
rect 19432 3392 19484 3398
rect 19432 3334 19484 3340
rect 19444 480 19472 3334
rect 20640 480 20668 3606
rect 21836 480 21864 7754
rect 22756 3466 22784 334562
rect 24214 3768 24270 3777
rect 23020 3732 23072 3738
rect 24214 3703 24270 3712
rect 23020 3674 23072 3680
rect 22744 3460 22796 3466
rect 22744 3402 22796 3408
rect 23032 480 23060 3674
rect 24228 480 24256 3703
rect 25320 3460 25372 3466
rect 25320 3402 25372 3408
rect 25332 480 25360 3402
rect 25516 3398 25544 336223
rect 35164 336048 35216 336054
rect 35164 335990 35216 335996
rect 29644 334688 29696 334694
rect 29644 334630 29696 334636
rect 26516 7880 26568 7886
rect 26516 7822 26568 7828
rect 25504 3392 25556 3398
rect 25504 3334 25556 3340
rect 26528 480 26556 7822
rect 28908 3596 28960 3602
rect 28908 3538 28960 3544
rect 27712 3052 27764 3058
rect 27712 2994 27764 3000
rect 27724 480 27752 2994
rect 28920 480 28948 3538
rect 29656 3058 29684 334630
rect 33784 331900 33836 331906
rect 33784 331842 33836 331848
rect 32404 329112 32456 329118
rect 32404 329054 32456 329060
rect 30104 7948 30156 7954
rect 30104 7890 30156 7896
rect 29644 3052 29696 3058
rect 29644 2994 29696 3000
rect 30116 480 30144 7890
rect 32416 6914 32444 329054
rect 33600 9036 33652 9042
rect 33600 8978 33652 8984
rect 32324 6886 32444 6914
rect 32324 3534 32352 6886
rect 32312 3528 32364 3534
rect 32312 3470 32364 3476
rect 32404 3528 32456 3534
rect 32404 3470 32456 3476
rect 31300 3392 31352 3398
rect 31300 3334 31352 3340
rect 31312 480 31340 3334
rect 32416 480 32444 3470
rect 33612 480 33640 8978
rect 33796 3398 33824 331842
rect 34796 4140 34848 4146
rect 34796 4082 34848 4088
rect 33784 3392 33836 3398
rect 33784 3334 33836 3340
rect 34808 480 34836 4082
rect 35176 3602 35204 335990
rect 39304 333260 39356 333266
rect 39304 333202 39356 333208
rect 36544 330540 36596 330546
rect 36544 330482 36596 330488
rect 36556 4146 36584 330482
rect 37188 9104 37240 9110
rect 37188 9046 37240 9052
rect 36544 4140 36596 4146
rect 36544 4082 36596 4088
rect 35992 3800 36044 3806
rect 35992 3742 36044 3748
rect 35164 3596 35216 3602
rect 35164 3538 35216 3544
rect 36004 480 36032 3742
rect 37200 480 37228 9046
rect 38384 3936 38436 3942
rect 38384 3878 38436 3884
rect 38396 480 38424 3878
rect 39316 3738 39344 333202
rect 41328 10328 41380 10334
rect 41328 10270 41380 10276
rect 39304 3732 39356 3738
rect 39304 3674 39356 3680
rect 39580 3664 39632 3670
rect 39580 3606 39632 3612
rect 39592 480 39620 3606
rect 41340 3602 41368 10270
rect 43076 4004 43128 4010
rect 43076 3946 43128 3952
rect 41880 3868 41932 3874
rect 41880 3810 41932 3816
rect 40684 3596 40736 3602
rect 40684 3538 40736 3544
rect 41328 3596 41380 3602
rect 41328 3538 41380 3544
rect 40696 480 40724 3538
rect 41892 480 41920 3810
rect 43088 480 43116 3946
rect 43456 3738 43484 336359
rect 114468 336330 114520 336336
rect 107568 336320 107620 336326
rect 107568 336262 107620 336268
rect 57244 336252 57296 336258
rect 57244 336194 57296 336200
rect 51724 336184 51776 336190
rect 51724 336126 51776 336132
rect 50344 336116 50396 336122
rect 50344 336058 50396 336064
rect 47584 329180 47636 329186
rect 47584 329122 47636 329128
rect 45468 10396 45520 10402
rect 45468 10338 45520 10344
rect 43444 3732 43496 3738
rect 43444 3674 43496 3680
rect 45376 3732 45428 3738
rect 45376 3674 45428 3680
rect 44272 3392 44324 3398
rect 44272 3334 44324 3340
rect 44284 480 44312 3334
rect 45388 1850 45416 3674
rect 45480 3398 45508 10338
rect 47596 3942 47624 329122
rect 49608 10464 49660 10470
rect 49608 10406 49660 10412
rect 47860 6180 47912 6186
rect 47860 6122 47912 6128
rect 47584 3936 47636 3942
rect 47584 3878 47636 3884
rect 45468 3392 45520 3398
rect 45468 3334 45520 3340
rect 46664 3392 46716 3398
rect 46664 3334 46716 3340
rect 45388 1822 45508 1850
rect 45480 480 45508 1822
rect 46676 480 46704 3334
rect 47872 480 47900 6122
rect 49620 3602 49648 10406
rect 50160 3936 50212 3942
rect 50160 3878 50212 3884
rect 48964 3596 49016 3602
rect 48964 3538 49016 3544
rect 49608 3596 49660 3602
rect 49608 3538 49660 3544
rect 48976 480 49004 3538
rect 50172 480 50200 3878
rect 50356 3806 50384 336058
rect 51356 6248 51408 6254
rect 51356 6190 51408 6196
rect 50344 3800 50396 3806
rect 50344 3742 50396 3748
rect 51368 480 51396 6190
rect 51736 4010 51764 336126
rect 54484 333328 54536 333334
rect 54484 333270 54536 333276
rect 53748 10532 53800 10538
rect 53748 10474 53800 10480
rect 51724 4004 51776 4010
rect 51724 3946 51776 3952
rect 53656 4004 53708 4010
rect 53656 3946 53708 3952
rect 52552 3596 52604 3602
rect 52552 3538 52604 3544
rect 52564 480 52592 3538
rect 53668 1986 53696 3946
rect 53760 3602 53788 10474
rect 54496 3874 54524 333270
rect 56508 10600 56560 10606
rect 56508 10542 56560 10548
rect 54944 6316 54996 6322
rect 54944 6258 54996 6264
rect 54484 3868 54536 3874
rect 54484 3810 54536 3816
rect 53748 3596 53800 3602
rect 53748 3538 53800 3544
rect 53668 1958 53788 1986
rect 53760 480 53788 1958
rect 54956 480 54984 6258
rect 56520 3398 56548 10542
rect 57256 4010 57284 336194
rect 87604 334824 87656 334830
rect 87604 334766 87656 334772
rect 86868 334756 86920 334762
rect 86868 334698 86920 334704
rect 84108 333396 84160 333402
rect 84108 333338 84160 333344
rect 68284 331968 68336 331974
rect 68284 331910 68336 331916
rect 58624 330608 58676 330614
rect 58624 330550 58676 330556
rect 58440 6384 58492 6390
rect 58440 6326 58492 6332
rect 57244 4004 57296 4010
rect 57244 3946 57296 3952
rect 56048 3392 56100 3398
rect 56048 3334 56100 3340
rect 56508 3392 56560 3398
rect 56508 3334 56560 3340
rect 56060 480 56088 3334
rect 57244 3188 57296 3194
rect 57244 3130 57296 3136
rect 57256 480 57284 3130
rect 58452 480 58480 6326
rect 58636 3738 58664 330550
rect 61384 329248 61436 329254
rect 61384 329190 61436 329196
rect 60648 10668 60700 10674
rect 60648 10610 60700 10616
rect 58624 3732 58676 3738
rect 58624 3674 58676 3680
rect 60660 3398 60688 10610
rect 60832 3732 60884 3738
rect 60832 3674 60884 3680
rect 59636 3392 59688 3398
rect 59636 3334 59688 3340
rect 60648 3392 60700 3398
rect 60648 3334 60700 3340
rect 59648 480 59676 3334
rect 60844 480 60872 3674
rect 61396 3194 61424 329190
rect 67548 10804 67600 10810
rect 67548 10746 67600 10752
rect 63224 10736 63276 10742
rect 63224 10678 63276 10684
rect 62028 6452 62080 6458
rect 62028 6394 62080 6400
rect 61384 3188 61436 3194
rect 61384 3130 61436 3136
rect 62040 480 62068 6394
rect 63236 480 63264 10678
rect 65524 6520 65576 6526
rect 65524 6462 65576 6468
rect 64328 3800 64380 3806
rect 64328 3742 64380 3748
rect 64340 480 64368 3742
rect 65536 480 65564 6462
rect 67560 3398 67588 10746
rect 68296 3942 68324 331910
rect 81348 330676 81400 330682
rect 81348 330618 81400 330624
rect 78588 11824 78640 11830
rect 78588 11766 78640 11772
rect 74448 11756 74500 11762
rect 74448 11698 74500 11704
rect 70308 10872 70360 10878
rect 70308 10814 70360 10820
rect 69112 6588 69164 6594
rect 69112 6530 69164 6536
rect 68284 3936 68336 3942
rect 68284 3878 68336 3884
rect 67916 3868 67968 3874
rect 67916 3810 67968 3816
rect 66720 3392 66772 3398
rect 66720 3334 66772 3340
rect 67548 3392 67600 3398
rect 67548 3334 67600 3340
rect 66732 480 66760 3334
rect 67928 480 67956 3810
rect 69124 480 69152 6530
rect 70320 480 70348 10814
rect 72608 8016 72660 8022
rect 72608 7958 72660 7964
rect 71504 3936 71556 3942
rect 71504 3878 71556 3884
rect 71516 480 71544 3878
rect 72620 480 72648 7958
rect 74460 3398 74488 11698
rect 76196 8084 76248 8090
rect 76196 8026 76248 8032
rect 75000 4004 75052 4010
rect 75000 3946 75052 3952
rect 73804 3392 73856 3398
rect 73804 3334 73856 3340
rect 74448 3392 74500 3398
rect 74448 3334 74500 3340
rect 73816 480 73844 3334
rect 75012 480 75040 3946
rect 76208 480 76236 8026
rect 78600 3398 78628 11766
rect 79692 8152 79744 8158
rect 79692 8094 79744 8100
rect 77392 3392 77444 3398
rect 77392 3334 77444 3340
rect 78588 3392 78640 3398
rect 78588 3334 78640 3340
rect 77404 480 77432 3334
rect 78588 3256 78640 3262
rect 78588 3198 78640 3204
rect 78600 480 78628 3198
rect 79704 480 79732 8094
rect 81360 3398 81388 330618
rect 82084 4072 82136 4078
rect 82084 4014 82136 4020
rect 80888 3392 80940 3398
rect 80888 3334 80940 3340
rect 81348 3392 81400 3398
rect 81348 3334 81400 3340
rect 80900 480 80928 3334
rect 82096 480 82124 4014
rect 84120 3330 84148 333338
rect 84476 3392 84528 3398
rect 84476 3334 84528 3340
rect 83280 3324 83332 3330
rect 83280 3266 83332 3272
rect 84108 3324 84160 3330
rect 84108 3266 84160 3272
rect 83292 480 83320 3266
rect 84488 480 84516 3334
rect 85672 3256 85724 3262
rect 85672 3198 85724 3204
rect 85684 480 85712 3198
rect 86880 480 86908 334698
rect 87616 3398 87644 334766
rect 93124 333532 93176 333538
rect 93124 333474 93176 333480
rect 88984 333464 89036 333470
rect 88984 333406 89036 333412
rect 87604 3392 87656 3398
rect 87604 3334 87656 3340
rect 88996 3330 89024 333406
rect 91008 10940 91060 10946
rect 91008 10882 91060 10888
rect 91020 3398 91048 10882
rect 93136 3398 93164 333474
rect 104164 332172 104216 332178
rect 104164 332114 104216 332120
rect 99288 332104 99340 332110
rect 99288 332046 99340 332052
rect 95148 332036 95200 332042
rect 95148 331978 95200 331984
rect 95056 11008 95108 11014
rect 95056 10950 95108 10956
rect 90364 3392 90416 3398
rect 90364 3334 90416 3340
rect 91008 3392 91060 3398
rect 91008 3334 91060 3340
rect 91560 3392 91612 3398
rect 91560 3334 91612 3340
rect 93124 3392 93176 3398
rect 93124 3334 93176 3340
rect 87972 3324 88024 3330
rect 87972 3266 88024 3272
rect 88984 3324 89036 3330
rect 88984 3266 89036 3272
rect 87984 480 88012 3266
rect 89168 3188 89220 3194
rect 89168 3130 89220 3136
rect 89180 480 89208 3130
rect 90376 480 90404 3334
rect 91572 480 91600 3334
rect 95068 3330 95096 10950
rect 93952 3324 94004 3330
rect 93952 3266 94004 3272
rect 95056 3324 95108 3330
rect 95056 3266 95108 3272
rect 92756 3256 92808 3262
rect 92756 3198 92808 3204
rect 92768 480 92796 3198
rect 93964 480 93992 3266
rect 95160 480 95188 331978
rect 97908 10260 97960 10266
rect 97908 10202 97960 10208
rect 97920 3330 97948 10202
rect 99300 3330 99328 332046
rect 102048 10192 102100 10198
rect 102048 10134 102100 10140
rect 102060 3330 102088 10134
rect 97448 3324 97500 3330
rect 97448 3266 97500 3272
rect 97908 3324 97960 3330
rect 97908 3266 97960 3272
rect 98644 3324 98696 3330
rect 98644 3266 98696 3272
rect 99288 3324 99340 3330
rect 99288 3266 99340 3272
rect 101036 3324 101088 3330
rect 101036 3266 101088 3272
rect 102048 3324 102100 3330
rect 102048 3266 102100 3272
rect 96252 3120 96304 3126
rect 96252 3062 96304 3068
rect 96264 480 96292 3062
rect 97460 480 97488 3266
rect 98656 480 98684 3266
rect 99840 2984 99892 2990
rect 99840 2926 99892 2932
rect 99852 480 99880 2926
rect 101048 480 101076 3266
rect 104176 3126 104204 332114
rect 106188 330744 106240 330750
rect 106188 330686 106240 330692
rect 104532 10124 104584 10130
rect 104532 10066 104584 10072
rect 102232 3120 102284 3126
rect 102232 3062 102284 3068
rect 104164 3120 104216 3126
rect 104164 3062 104216 3068
rect 102244 480 102272 3062
rect 103336 3052 103388 3058
rect 103336 2994 103388 3000
rect 103348 480 103376 2994
rect 104544 480 104572 10066
rect 106200 3126 106228 330686
rect 107580 3126 107608 336262
rect 111064 330812 111116 330818
rect 111064 330754 111116 330760
rect 108948 10056 109000 10062
rect 108948 9998 109000 10004
rect 108960 3126 108988 9998
rect 111076 3126 111104 330754
rect 113088 329316 113140 329322
rect 113088 329258 113140 329264
rect 111616 9988 111668 9994
rect 111616 9930 111668 9936
rect 105728 3120 105780 3126
rect 105728 3062 105780 3068
rect 106188 3120 106240 3126
rect 106188 3062 106240 3068
rect 106924 3120 106976 3126
rect 106924 3062 106976 3068
rect 107568 3120 107620 3126
rect 107568 3062 107620 3068
rect 108120 3120 108172 3126
rect 108120 3062 108172 3068
rect 108948 3120 109000 3126
rect 108948 3062 109000 3068
rect 109316 3120 109368 3126
rect 109316 3062 109368 3068
rect 111064 3120 111116 3126
rect 111064 3062 111116 3068
rect 105740 480 105768 3062
rect 106936 480 106964 3062
rect 108132 480 108160 3062
rect 109328 480 109356 3062
rect 110512 2984 110564 2990
rect 110512 2926 110564 2932
rect 110524 480 110552 2926
rect 111628 480 111656 9930
rect 113100 6914 113128 329258
rect 112824 6886 113128 6914
rect 112824 480 112852 6886
rect 114480 2922 114508 336330
rect 117228 330880 117280 330886
rect 117228 330822 117280 330828
rect 115848 9920 115900 9926
rect 115848 9862 115900 9868
rect 115860 2922 115888 9862
rect 117240 2922 117268 330822
rect 124128 329452 124180 329458
rect 124128 329394 124180 329400
rect 119988 329384 120040 329390
rect 119988 329326 120040 329332
rect 119804 9852 119856 9858
rect 119804 9794 119856 9800
rect 119816 2922 119844 9794
rect 120000 6914 120028 329326
rect 122748 9784 122800 9790
rect 122748 9726 122800 9732
rect 119908 6886 120028 6914
rect 114008 2916 114060 2922
rect 114008 2858 114060 2864
rect 114468 2916 114520 2922
rect 114468 2858 114520 2864
rect 115204 2916 115256 2922
rect 115204 2858 115256 2864
rect 115848 2916 115900 2922
rect 115848 2858 115900 2864
rect 116400 2916 116452 2922
rect 116400 2858 116452 2864
rect 117228 2916 117280 2922
rect 117228 2858 117280 2864
rect 118792 2916 118844 2922
rect 118792 2858 118844 2864
rect 119804 2916 119856 2922
rect 119804 2858 119856 2864
rect 114020 480 114048 2858
rect 115216 480 115244 2858
rect 116412 480 116440 2858
rect 117596 2848 117648 2854
rect 117596 2790 117648 2796
rect 117608 480 117636 2790
rect 118804 480 118832 2858
rect 119908 480 119936 6886
rect 122760 2922 122788 9726
rect 124140 2922 124168 329394
rect 125520 6914 125548 336398
rect 204904 335980 204956 335986
rect 204904 335922 204956 335928
rect 197268 335300 197320 335306
rect 197268 335242 197320 335248
rect 179328 335232 179380 335238
rect 179328 335174 179380 335180
rect 169668 335164 169720 335170
rect 169668 335106 169720 335112
rect 161388 335096 161440 335102
rect 161388 335038 161440 335044
rect 144828 335028 144880 335034
rect 144828 334970 144880 334976
rect 140688 334892 140740 334898
rect 140688 334834 140740 334840
rect 138848 15904 138900 15910
rect 138848 15846 138900 15852
rect 125876 13320 125928 13326
rect 125876 13262 125928 13268
rect 125428 6886 125548 6914
rect 125428 2922 125456 6886
rect 122288 2916 122340 2922
rect 122288 2858 122340 2864
rect 122748 2916 122800 2922
rect 122748 2858 122800 2864
rect 123484 2916 123536 2922
rect 123484 2858 123536 2864
rect 124128 2916 124180 2922
rect 124128 2858 124180 2864
rect 124680 2916 124732 2922
rect 124680 2858 124732 2864
rect 125416 2916 125468 2922
rect 125416 2858 125468 2864
rect 121092 2848 121144 2854
rect 121092 2790 121144 2796
rect 121104 480 121132 2790
rect 122300 480 122328 2858
rect 123496 480 123524 2858
rect 124692 480 124720 2858
rect 125888 480 125916 13262
rect 128176 13116 128228 13122
rect 128176 13058 128228 13064
rect 126980 8900 127032 8906
rect 126980 8842 127032 8848
rect 126992 480 127020 8842
rect 128188 480 128216 13058
rect 135260 9240 135312 9246
rect 135260 9182 135312 9188
rect 131764 9172 131816 9178
rect 131764 9114 131816 9120
rect 130568 6656 130620 6662
rect 130568 6598 130620 6604
rect 129372 5092 129424 5098
rect 129372 5034 129424 5040
rect 129384 480 129412 5034
rect 130580 480 130608 6598
rect 131776 480 131804 9114
rect 134156 8220 134208 8226
rect 134156 8162 134208 8168
rect 132960 5160 133012 5166
rect 132960 5102 133012 5108
rect 132972 480 133000 5102
rect 134168 480 134196 8162
rect 135272 480 135300 9182
rect 137652 8288 137704 8294
rect 137652 8230 137704 8236
rect 136456 5296 136508 5302
rect 136456 5238 136508 5244
rect 136468 480 136496 5238
rect 137664 480 137692 8230
rect 138860 480 138888 15846
rect 140700 6914 140728 334834
rect 143448 332240 143500 332246
rect 143448 332182 143500 332188
rect 141240 7540 141292 7546
rect 141240 7482 141292 7488
rect 140056 6886 140728 6914
rect 140056 480 140084 6886
rect 141252 480 141280 7482
rect 143460 6914 143488 332182
rect 144736 7472 144788 7478
rect 144736 7414 144788 7420
rect 142448 6886 143488 6914
rect 142448 480 142476 6886
rect 143540 4208 143592 4214
rect 143540 4150 143592 4156
rect 143552 480 143580 4150
rect 144748 480 144776 7414
rect 144840 4214 144868 334970
rect 147588 334960 147640 334966
rect 147588 334902 147640 334908
rect 146208 330948 146260 330954
rect 146208 330890 146260 330896
rect 146220 6914 146248 330890
rect 147600 6914 147628 334902
rect 158628 333668 158680 333674
rect 158628 333610 158680 333616
rect 151728 333600 151780 333606
rect 151728 333542 151780 333548
rect 149520 13184 149572 13190
rect 149520 13126 149572 13132
rect 148324 7404 148376 7410
rect 148324 7346 148376 7352
rect 145944 6886 146248 6914
rect 147140 6886 147628 6914
rect 144828 4208 144880 4214
rect 144828 4150 144880 4156
rect 145944 480 145972 6886
rect 147140 480 147168 6886
rect 148336 480 148364 7346
rect 149532 480 149560 13126
rect 151740 6914 151768 333542
rect 153108 331016 153160 331022
rect 153108 330958 153160 330964
rect 151820 7336 151872 7342
rect 151820 7278 151872 7284
rect 150636 6886 151768 6914
rect 150636 480 150664 6886
rect 151832 480 151860 7278
rect 153120 6914 153148 330958
rect 157248 18624 157300 18630
rect 157248 18566 157300 18572
rect 154212 11960 154264 11966
rect 154212 11902 154264 11908
rect 153028 6886 153148 6914
rect 153028 480 153056 6886
rect 154224 480 154252 11902
rect 155408 7268 155460 7274
rect 155408 7210 155460 7216
rect 155420 480 155448 7210
rect 157260 6914 157288 18566
rect 158640 6914 158668 333610
rect 161296 17264 161348 17270
rect 161296 17206 161348 17212
rect 161308 11694 161336 17206
rect 160100 11688 160152 11694
rect 160100 11630 160152 11636
rect 161296 11688 161348 11694
rect 161296 11630 161348 11636
rect 158904 7200 158956 7206
rect 158904 7142 158956 7148
rect 156616 6886 157288 6914
rect 157812 6886 158668 6914
rect 156616 480 156644 6886
rect 157812 480 157840 6886
rect 158916 480 158944 7142
rect 160112 480 160140 11630
rect 161400 6914 161428 335038
rect 162768 333736 162820 333742
rect 162768 333678 162820 333684
rect 162780 6914 162808 333678
rect 163688 13252 163740 13258
rect 163688 13194 163740 13200
rect 161308 6886 161428 6914
rect 162504 6886 162808 6914
rect 161308 480 161336 6886
rect 162504 480 162532 6886
rect 163700 480 163728 13194
rect 164884 12028 164936 12034
rect 164884 11970 164936 11976
rect 164896 480 164924 11970
rect 167184 11892 167236 11898
rect 167184 11834 167236 11840
rect 166080 6724 166132 6730
rect 166080 6666 166132 6672
rect 166092 480 166120 6666
rect 167196 480 167224 11834
rect 169576 6792 169628 6798
rect 169576 6734 169628 6740
rect 168380 1692 168432 1698
rect 168380 1634 168432 1640
rect 168392 480 168420 1634
rect 169588 480 169616 6734
rect 169680 1698 169708 335106
rect 177948 333804 178000 333810
rect 177948 333746 178000 333752
rect 175188 332376 175240 332382
rect 175188 332318 175240 332324
rect 171048 332308 171100 332314
rect 171048 332250 171100 332256
rect 171060 6914 171088 332250
rect 175200 6914 175228 332318
rect 175464 12096 175516 12102
rect 175464 12038 175516 12044
rect 170784 6886 171088 6914
rect 174280 6886 175228 6914
rect 169668 1692 169720 1698
rect 169668 1634 169720 1640
rect 170784 480 170812 6886
rect 173164 6112 173216 6118
rect 173164 6054 173216 6060
rect 171968 4684 172020 4690
rect 171968 4626 172020 4632
rect 171980 480 172008 4626
rect 173176 480 173204 6054
rect 174280 480 174308 6886
rect 175476 480 175504 12038
rect 177960 6914 177988 333746
rect 179340 6914 179368 335174
rect 188988 332512 189040 332518
rect 188988 332454 189040 332460
rect 182088 332444 182140 332450
rect 182088 332386 182140 332392
rect 182100 6914 182128 332386
rect 186136 13388 186188 13394
rect 186136 13330 186188 13336
rect 182548 12164 182600 12170
rect 182548 12106 182600 12112
rect 177868 6886 177988 6914
rect 179064 6886 179368 6914
rect 181456 6886 182128 6914
rect 176660 6044 176712 6050
rect 176660 5986 176712 5992
rect 176672 480 176700 5986
rect 177868 480 177896 6886
rect 179064 480 179092 6886
rect 180248 5976 180300 5982
rect 180248 5918 180300 5924
rect 180260 480 180288 5918
rect 181456 480 181484 6886
rect 182560 480 182588 12106
rect 183744 5908 183796 5914
rect 183744 5850 183796 5856
rect 183756 480 183784 5850
rect 186148 4214 186176 13330
rect 189000 6914 189028 332454
rect 195612 9376 195664 9382
rect 195612 9318 195664 9324
rect 192024 9308 192076 9314
rect 192024 9250 192076 9256
rect 188540 6886 189028 6914
rect 187332 5840 187384 5846
rect 187332 5782 187384 5788
rect 186228 5500 186280 5506
rect 186228 5442 186280 5448
rect 184940 4208 184992 4214
rect 184940 4150 184992 4156
rect 186136 4208 186188 4214
rect 186136 4150 186188 4156
rect 184952 480 184980 4150
rect 186240 2802 186268 5442
rect 186148 2774 186268 2802
rect 186148 480 186176 2774
rect 187344 480 187372 5782
rect 188540 480 188568 6886
rect 190828 5772 190880 5778
rect 190828 5714 190880 5720
rect 189724 5432 189776 5438
rect 189724 5374 189776 5380
rect 189736 480 189764 5374
rect 190840 480 190868 5714
rect 192036 480 192064 9250
rect 194416 5704 194468 5710
rect 194416 5646 194468 5652
rect 193220 4752 193272 4758
rect 193220 4694 193272 4700
rect 193232 480 193260 4694
rect 194428 480 194456 5646
rect 195624 480 195652 9318
rect 197280 6914 197308 335242
rect 202788 334552 202840 334558
rect 202788 334494 202840 334500
rect 198648 333872 198700 333878
rect 198648 333814 198700 333820
rect 198660 6914 198688 333814
rect 202696 9512 202748 9518
rect 202696 9454 202748 9460
rect 199108 9444 199160 9450
rect 199108 9386 199160 9392
rect 196820 6886 197308 6914
rect 197924 6886 198688 6914
rect 196820 480 196848 6886
rect 197924 480 197952 6886
rect 199120 480 199148 9386
rect 200304 4276 200356 4282
rect 200304 4218 200356 4224
rect 200316 480 200344 4218
rect 201500 4208 201552 4214
rect 201500 4150 201552 4156
rect 201512 480 201540 4150
rect 202708 480 202736 9454
rect 202800 4214 202828 334494
rect 204916 5302 204944 335922
rect 205548 333940 205600 333946
rect 205548 333882 205600 333888
rect 205560 6914 205588 333882
rect 209056 16574 209084 336466
rect 213184 335640 213236 335646
rect 213184 335582 213236 335588
rect 209688 333192 209740 333198
rect 209688 333134 209740 333140
rect 208964 16546 209084 16574
rect 206192 9580 206244 9586
rect 206192 9522 206244 9528
rect 205100 6886 205588 6914
rect 204904 5296 204956 5302
rect 204904 5238 204956 5244
rect 203892 5228 203944 5234
rect 203892 5170 203944 5176
rect 202788 4208 202840 4214
rect 202788 4150 202840 4156
rect 203904 480 203932 5170
rect 205100 480 205128 6886
rect 206204 480 206232 9522
rect 207388 5296 207440 5302
rect 207388 5238 207440 5244
rect 207400 480 207428 5238
rect 208964 4282 208992 16546
rect 209700 6914 209728 333134
rect 212172 12232 212224 12238
rect 212172 12174 212224 12180
rect 209780 9648 209832 9654
rect 209780 9590 209832 9596
rect 209056 6886 209728 6914
rect 208952 4276 209004 4282
rect 208952 4218 209004 4224
rect 209056 3482 209084 6886
rect 208596 3454 209084 3482
rect 208596 480 208624 3454
rect 209792 480 209820 9590
rect 210976 5364 211028 5370
rect 210976 5306 211028 5312
rect 210988 480 211016 5306
rect 212184 480 212212 12174
rect 213196 8906 213224 335582
rect 213184 8900 213236 8906
rect 213184 8842 213236 8848
rect 213368 8900 213420 8906
rect 213368 8842 213420 8848
rect 213380 480 213408 8842
rect 214576 6914 214604 336534
rect 214300 6886 214604 6914
rect 214300 5438 214328 6886
rect 215956 5506 215984 336602
rect 216588 334484 216640 334490
rect 216588 334426 216640 334432
rect 216600 6914 216628 334426
rect 219256 332580 219308 332586
rect 219256 332522 219308 332528
rect 216864 8832 216916 8838
rect 216864 8774 216916 8780
rect 216048 6886 216628 6914
rect 215944 5500 215996 5506
rect 215944 5442 215996 5448
rect 214288 5432 214340 5438
rect 214288 5374 214340 5380
rect 214472 5432 214524 5438
rect 214472 5374 214524 5380
rect 214484 480 214512 5374
rect 216048 3482 216076 6886
rect 215680 3454 216076 3482
rect 215680 480 215708 3454
rect 216876 480 216904 8774
rect 218060 5500 218112 5506
rect 218060 5442 218112 5448
rect 218072 480 218100 5442
rect 219268 480 219296 332522
rect 220096 4758 220124 336670
rect 224224 335912 224276 335918
rect 224224 335854 224276 335860
rect 222844 335776 222896 335782
rect 222844 335718 222896 335724
rect 220452 8764 220504 8770
rect 220452 8706 220504 8712
rect 220084 4752 220136 4758
rect 220084 4694 220136 4700
rect 220464 480 220492 8706
rect 221556 4752 221608 4758
rect 221556 4694 221608 4700
rect 221568 480 221596 4694
rect 222856 4690 222884 335718
rect 223488 334416 223540 334422
rect 223488 334358 223540 334364
rect 223500 6914 223528 334358
rect 224236 12170 224264 335854
rect 226984 335708 227036 335714
rect 226984 335650 227036 335656
rect 224224 12164 224276 12170
rect 224224 12106 224276 12112
rect 226996 12102 227024 335650
rect 227628 333124 227680 333130
rect 227628 333066 227680 333072
rect 226984 12096 227036 12102
rect 226984 12038 227036 12044
rect 223948 8696 224000 8702
rect 223948 8638 224000 8644
rect 222948 6886 223528 6914
rect 222844 4684 222896 4690
rect 222844 4626 222896 4632
rect 222948 3482 222976 6886
rect 222764 3454 222976 3482
rect 222764 480 222792 3454
rect 223960 480 223988 8638
rect 227536 8628 227588 8634
rect 227536 8570 227588 8576
rect 225144 4684 225196 4690
rect 225144 4626 225196 4632
rect 225156 480 225184 4626
rect 226340 4208 226392 4214
rect 226340 4150 226392 4156
rect 226352 480 226380 4150
rect 227548 480 227576 8570
rect 227640 4214 227668 333066
rect 228376 45558 228404 458322
rect 231136 398818 231164 458730
rect 232596 458516 232648 458522
rect 232596 458458 232648 458464
rect 231124 398812 231176 398818
rect 231124 398754 231176 398760
rect 231124 335572 231176 335578
rect 231124 335514 231176 335520
rect 228364 45552 228416 45558
rect 228364 45494 228416 45500
rect 231136 12034 231164 335514
rect 232504 335504 232556 335510
rect 232504 335446 232556 335452
rect 231124 12028 231176 12034
rect 231124 11970 231176 11976
rect 232516 11966 232544 335446
rect 232608 215286 232636 458458
rect 267476 457994 267504 459546
rect 270408 458448 270460 458454
rect 270408 458390 270460 458396
rect 269028 458312 269080 458318
rect 269028 458254 269080 458260
rect 269040 457994 269068 458254
rect 267352 457966 267504 457994
rect 268916 457966 269068 457994
rect 270420 457994 270448 458390
rect 272352 457994 272380 459614
rect 273996 458856 274048 458862
rect 273996 458798 274048 458804
rect 274008 457994 274036 458798
rect 280068 458720 280120 458726
rect 280068 458662 280120 458668
rect 277032 458584 277084 458590
rect 277032 458526 277084 458532
rect 277044 457994 277072 458526
rect 280080 457994 280108 458662
rect 270420 457966 270480 457994
rect 272044 457966 272380 457994
rect 273700 457966 274036 457994
rect 276828 457966 277072 457994
rect 279956 457966 280108 457994
rect 281460 457994 281488 459750
rect 285600 459746 285628 484366
rect 286968 470620 287020 470626
rect 286968 470562 287020 470568
rect 286980 460934 287008 470562
rect 288360 460934 288388 510614
rect 286704 460906 287008 460934
rect 288268 460906 288388 460934
rect 285036 459740 285088 459746
rect 285036 459682 285088 459688
rect 285588 459740 285640 459746
rect 285588 459682 285640 459688
rect 285048 457994 285076 459682
rect 286704 457994 286732 460906
rect 288268 457994 288296 460906
rect 289740 457994 289768 536794
rect 291108 524476 291160 524482
rect 291108 524418 291160 524424
rect 291120 457994 291148 524418
rect 293880 459814 293908 563042
rect 295260 459814 295288 590650
rect 296628 576904 296680 576910
rect 296628 576846 296680 576852
rect 296640 459814 296668 576846
rect 298020 460934 298048 616830
rect 299400 460934 299428 643078
rect 300676 630692 300728 630698
rect 300676 630634 300728 630640
rect 297744 460906 298048 460934
rect 299308 460906 299428 460934
rect 292948 459808 293000 459814
rect 292948 459750 293000 459756
rect 293868 459808 293920 459814
rect 293868 459750 293920 459756
rect 294512 459808 294564 459814
rect 294512 459750 294564 459756
rect 295248 459808 295300 459814
rect 295248 459750 295300 459756
rect 296076 459808 296128 459814
rect 296076 459750 296128 459756
rect 296628 459808 296680 459814
rect 296628 459750 296680 459756
rect 292960 457994 292988 459750
rect 294524 457994 294552 459750
rect 296088 457994 296116 459750
rect 297744 457994 297772 460906
rect 299308 457994 299336 460906
rect 300688 457994 300716 630634
rect 300780 459882 300808 699654
rect 304908 696992 304960 696998
rect 304908 696934 304960 696940
rect 302148 670812 302200 670818
rect 302148 670754 302200 670760
rect 300768 459876 300820 459882
rect 300768 459818 300820 459824
rect 302160 458266 302188 670754
rect 304920 459814 304948 696934
rect 306288 683188 306340 683194
rect 306288 683130 306340 683136
rect 306300 459814 306328 683130
rect 307680 459814 307708 700402
rect 309060 460934 309088 700538
rect 310428 700528 310480 700534
rect 310428 700470 310480 700476
rect 310440 460934 310468 700470
rect 308784 460906 309088 460934
rect 310348 460906 310468 460934
rect 303988 459808 304040 459814
rect 303988 459750 304040 459756
rect 304908 459808 304960 459814
rect 304908 459750 304960 459756
rect 305552 459808 305604 459814
rect 305552 459750 305604 459756
rect 306288 459808 306340 459814
rect 306288 459750 306340 459756
rect 307116 459808 307168 459814
rect 307116 459750 307168 459756
rect 307668 459808 307720 459814
rect 307668 459750 307720 459756
rect 281460 457966 281520 457994
rect 284740 457966 285076 457994
rect 286304 457966 286732 457994
rect 287868 457966 288296 457994
rect 289432 457966 289768 457994
rect 290996 457966 291148 457994
rect 292652 457966 292988 457994
rect 294216 457966 294552 457994
rect 295780 457966 296116 457994
rect 297344 457966 297772 457994
rect 298908 457966 299336 457994
rect 300472 457966 300716 457994
rect 302114 458238 302188 458266
rect 302114 457980 302142 458238
rect 304000 457994 304028 459750
rect 305564 457994 305592 459750
rect 307128 457994 307156 459750
rect 308784 457994 308812 460906
rect 310348 457994 310376 460906
rect 311820 457994 311848 700674
rect 313200 458266 313228 700810
rect 315948 700800 316000 700806
rect 315948 700742 316000 700748
rect 315960 459814 315988 700742
rect 317340 459814 317368 700946
rect 331312 700936 331364 700942
rect 331312 700878 331364 700884
rect 320088 700256 320140 700262
rect 320088 700198 320140 700204
rect 318708 700188 318760 700194
rect 318708 700130 318760 700136
rect 318720 459814 318748 700130
rect 320100 460934 320128 700198
rect 327080 700120 327132 700126
rect 327080 700062 327132 700068
rect 321468 700052 321520 700058
rect 321468 699994 321520 700000
rect 319824 460906 320128 460934
rect 315028 459808 315080 459814
rect 315028 459750 315080 459756
rect 315948 459808 316000 459814
rect 315948 459750 316000 459756
rect 316592 459808 316644 459814
rect 316592 459750 316644 459756
rect 317328 459808 317380 459814
rect 317328 459750 317380 459756
rect 318156 459808 318208 459814
rect 318156 459750 318208 459756
rect 318708 459808 318760 459814
rect 318708 459750 318760 459756
rect 303692 457966 304028 457994
rect 305256 457966 305592 457994
rect 306820 457966 307156 457994
rect 308384 457966 308812 457994
rect 309948 457966 310376 457994
rect 311604 457966 311848 457994
rect 313154 458238 313228 458266
rect 313154 457980 313182 458238
rect 315040 457994 315068 459750
rect 316604 457994 316632 459750
rect 318168 457994 318196 459750
rect 319824 457994 319852 460906
rect 321480 457994 321508 699994
rect 324228 699984 324280 699990
rect 324228 699926 324280 699932
rect 322848 699916 322900 699922
rect 322848 699858 322900 699864
rect 322860 457994 322888 699858
rect 324240 458266 324268 699926
rect 325700 459944 325752 459950
rect 325700 459886 325752 459892
rect 314732 457966 315068 457994
rect 316296 457966 316632 457994
rect 317860 457966 318196 457994
rect 319424 457966 319852 457994
rect 321080 457966 321508 457994
rect 322644 457966 322888 457994
rect 324194 458238 324268 458266
rect 324194 457980 324222 458238
rect 325712 457994 325740 459886
rect 327092 457994 327120 700062
rect 331324 480254 331352 700878
rect 332520 699922 332548 703520
rect 336740 700664 336792 700670
rect 336740 700606 336792 700612
rect 332508 699916 332560 699922
rect 332508 699858 332560 699864
rect 333244 670744 333296 670750
rect 333244 670686 333296 670692
rect 331324 480226 331720 480254
rect 330208 460080 330260 460086
rect 330208 460022 330260 460028
rect 328552 460012 328604 460018
rect 328552 459954 328604 459960
rect 328564 457994 328592 459954
rect 330220 457994 330248 460022
rect 331692 457994 331720 480226
rect 333256 460154 333284 670686
rect 334900 460896 334952 460902
rect 334900 460838 334952 460844
rect 333244 460148 333296 460154
rect 333244 460090 333296 460096
rect 333336 460080 333388 460086
rect 333336 460022 333388 460028
rect 333348 457994 333376 460022
rect 334912 457994 334940 460838
rect 336752 457994 336780 700606
rect 340880 700392 340932 700398
rect 340880 700334 340932 700340
rect 338764 618316 338816 618322
rect 338764 618258 338816 618264
rect 338776 460834 338804 618258
rect 340892 480254 340920 700334
rect 345020 700324 345072 700330
rect 345020 700266 345072 700272
rect 342904 565888 342956 565894
rect 342904 565830 342956 565836
rect 340892 480226 341196 480254
rect 338120 460828 338172 460834
rect 338120 460770 338172 460776
rect 338764 460828 338816 460834
rect 338764 460770 338816 460776
rect 338132 457994 338160 460770
rect 339684 460760 339736 460766
rect 339684 460702 339736 460708
rect 339696 457994 339724 460702
rect 341168 457994 341196 480226
rect 342916 460698 342944 565830
rect 345032 480254 345060 700266
rect 348804 699990 348832 703520
rect 364996 700058 365024 703520
rect 397472 700194 397500 703520
rect 413664 700262 413692 703520
rect 429856 701010 429884 703520
rect 429844 701004 429896 701010
rect 429844 700946 429896 700952
rect 462332 700874 462360 703520
rect 462320 700868 462372 700874
rect 462320 700810 462372 700816
rect 478524 700806 478552 703520
rect 478512 700800 478564 700806
rect 478512 700742 478564 700748
rect 494808 700738 494836 703520
rect 494796 700732 494848 700738
rect 494796 700674 494848 700680
rect 527192 700602 527220 703520
rect 527180 700596 527232 700602
rect 527180 700538 527232 700544
rect 543476 700534 543504 703520
rect 543464 700528 543516 700534
rect 543464 700470 543516 700476
rect 559668 700466 559696 703520
rect 559656 700460 559708 700466
rect 559656 700402 559708 700408
rect 413652 700256 413704 700262
rect 413652 700198 413704 700204
rect 397460 700188 397512 700194
rect 397460 700130 397512 700136
rect 364984 700052 365036 700058
rect 364984 699994 365036 700000
rect 348792 699984 348844 699990
rect 348792 699926 348844 699932
rect 580170 697232 580226 697241
rect 580170 697167 580226 697176
rect 580184 696998 580212 697167
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 580170 683904 580226 683913
rect 580170 683839 580226 683848
rect 580184 683194 580212 683839
rect 580172 683188 580224 683194
rect 580172 683130 580224 683136
rect 580172 670812 580224 670818
rect 580172 670754 580224 670760
rect 580184 670721 580212 670754
rect 580170 670712 580226 670721
rect 580170 670647 580226 670656
rect 350540 656940 350592 656946
rect 350540 656882 350592 656888
rect 348424 514820 348476 514826
rect 348424 514762 348476 514768
rect 345032 480226 345888 480254
rect 342812 460692 342864 460698
rect 342812 460634 342864 460640
rect 342904 460692 342956 460698
rect 342904 460634 342956 460640
rect 342824 457994 342852 460634
rect 344376 460624 344428 460630
rect 344376 460566 344428 460572
rect 344388 457994 344416 460566
rect 345860 457994 345888 480226
rect 348436 460562 348464 514762
rect 350552 480254 350580 656882
rect 580170 644056 580226 644065
rect 580170 643991 580226 644000
rect 580184 643142 580212 643991
rect 580172 643136 580224 643142
rect 580172 643078 580224 643084
rect 580170 630864 580226 630873
rect 580170 630799 580226 630808
rect 580184 630698 580212 630799
rect 580172 630692 580224 630698
rect 580172 630634 580224 630640
rect 580170 617536 580226 617545
rect 580170 617471 580226 617480
rect 580184 616894 580212 617471
rect 580172 616888 580224 616894
rect 580172 616830 580224 616836
rect 354680 605872 354732 605878
rect 354680 605814 354732 605820
rect 354692 480254 354720 605814
rect 579802 591016 579858 591025
rect 579802 590951 579858 590960
rect 579816 590714 579844 590951
rect 579804 590708 579856 590714
rect 579804 590650 579856 590656
rect 580170 577688 580226 577697
rect 580170 577623 580226 577632
rect 580184 576910 580212 577623
rect 580172 576904 580224 576910
rect 580172 576846 580224 576852
rect 579802 564360 579858 564369
rect 579802 564295 579858 564304
rect 579816 563106 579844 564295
rect 579804 563100 579856 563106
rect 579804 563042 579856 563048
rect 360200 553444 360252 553450
rect 360200 553386 360252 553392
rect 350552 480226 350672 480254
rect 354692 480226 355364 480254
rect 347780 460556 347832 460562
rect 347780 460498 347832 460504
rect 348424 460556 348476 460562
rect 348424 460498 348476 460504
rect 347792 457994 347820 460498
rect 349160 460488 349212 460494
rect 349160 460430 349212 460436
rect 349172 457994 349200 460430
rect 350644 457994 350672 480226
rect 352564 462392 352616 462398
rect 352564 462334 352616 462340
rect 352576 460494 352604 462334
rect 352564 460488 352616 460494
rect 352564 460430 352616 460436
rect 353852 460420 353904 460426
rect 353852 460362 353904 460368
rect 352288 460148 352340 460154
rect 352288 460090 352340 460096
rect 352300 457994 352328 460090
rect 353864 457994 353892 460362
rect 355336 457994 355364 480226
rect 356980 460828 357032 460834
rect 356980 460770 357032 460776
rect 356992 457994 357020 460770
rect 358820 460352 358872 460358
rect 358820 460294 358872 460300
rect 358832 457994 358860 460294
rect 360212 457994 360240 553386
rect 580170 537840 580226 537849
rect 580170 537775 580226 537784
rect 580184 536858 580212 537775
rect 580172 536852 580224 536858
rect 580172 536794 580224 536800
rect 580170 524512 580226 524521
rect 580170 524447 580172 524456
rect 580224 524447 580226 524456
rect 580172 524418 580224 524424
rect 580170 511320 580226 511329
rect 580170 511255 580226 511264
rect 580184 510678 580212 511255
rect 580172 510672 580224 510678
rect 580172 510614 580224 510620
rect 364340 501016 364392 501022
rect 364340 500958 364392 500964
rect 364352 480254 364380 500958
rect 580170 484664 580226 484673
rect 580170 484599 580226 484608
rect 580184 484430 580212 484599
rect 580172 484424 580224 484430
rect 580172 484366 580224 484372
rect 364352 480226 364840 480254
rect 361764 460692 361816 460698
rect 361764 460634 361816 460640
rect 361776 457994 361804 460634
rect 363328 460284 363380 460290
rect 363328 460226 363380 460232
rect 363340 457994 363368 460226
rect 364812 457994 364840 480226
rect 579986 471472 580042 471481
rect 579986 471407 580042 471416
rect 580000 470626 580028 471407
rect 579988 470620 580040 470626
rect 579988 470562 580040 470568
rect 366456 460556 366508 460562
rect 366456 460498 366508 460504
rect 366468 457994 366496 460498
rect 371240 460488 371292 460494
rect 371240 460430 371292 460436
rect 368112 460216 368164 460222
rect 368112 460158 368164 460164
rect 368124 457994 368152 460158
rect 371252 457994 371280 460430
rect 569224 459740 569276 459746
rect 569224 459682 569276 459688
rect 566464 459672 566516 459678
rect 566464 459614 566516 459620
rect 562324 459604 562376 459610
rect 562324 459546 562376 459552
rect 416044 458856 416096 458862
rect 416044 458798 416096 458804
rect 374368 458788 374420 458794
rect 374368 458730 374420 458736
rect 373126 458244 373178 458250
rect 373126 458186 373178 458192
rect 325712 457966 325772 457994
rect 327092 457966 327336 457994
rect 328564 457966 328900 457994
rect 330220 457966 330556 457994
rect 331692 457966 332120 457994
rect 333348 457966 333684 457994
rect 334912 457966 335248 457994
rect 336752 457966 336812 457994
rect 338132 457966 338376 457994
rect 339696 457966 340032 457994
rect 341168 457966 341596 457994
rect 342824 457966 343160 457994
rect 344388 457966 344724 457994
rect 345860 457966 346288 457994
rect 347792 457966 347852 457994
rect 349172 457966 349508 457994
rect 350644 457966 351072 457994
rect 352300 457966 352636 457994
rect 353864 457966 354200 457994
rect 355336 457966 355764 457994
rect 356992 457966 357328 457994
rect 358832 457966 358984 457994
rect 360212 457966 360548 457994
rect 361776 457966 362112 457994
rect 363340 457966 363676 457994
rect 364812 457966 365240 457994
rect 366468 457966 366804 457994
rect 368124 457966 368460 457994
rect 371252 457966 371588 457994
rect 373138 457980 373166 458186
rect 374380 457994 374408 458730
rect 375932 458652 375984 458658
rect 375932 458594 375984 458600
rect 375944 457994 375972 458594
rect 391940 458516 391992 458522
rect 391940 458458 391992 458464
rect 391952 457994 391980 458458
rect 407580 458380 407632 458386
rect 407580 458322 407632 458328
rect 407592 457994 407620 458322
rect 374380 457966 374716 457994
rect 375944 457966 376280 457994
rect 391952 457966 392104 457994
rect 407592 457966 407928 457994
rect 283472 457496 283524 457502
rect 283176 457444 283472 457450
rect 283176 457438 283524 457444
rect 233884 457428 233936 457434
rect 283176 457422 283512 457438
rect 369872 457434 370024 457450
rect 377600 457434 377936 457450
rect 379164 457434 379500 457450
rect 380912 457434 381064 457450
rect 369860 457428 370024 457434
rect 233884 457370 233936 457376
rect 369912 457422 370024 457428
rect 377588 457428 377936 457434
rect 369860 457370 369912 457376
rect 377640 457422 377936 457428
rect 379152 457428 379500 457434
rect 377588 457370 377640 457376
rect 379204 457422 379500 457428
rect 380900 457428 381064 457434
rect 379152 457370 379204 457376
rect 380952 457422 381064 457428
rect 380900 457370 380952 457376
rect 233896 449886 233924 457370
rect 278688 457360 278740 457366
rect 237194 457328 237250 457337
rect 234632 457286 235796 457314
rect 233884 449880 233936 449886
rect 233884 449822 233936 449828
rect 233884 335844 233936 335850
rect 233884 335786 233936 335792
rect 232596 215280 232648 215286
rect 232596 215222 232648 215228
rect 233896 12238 233924 335786
rect 233976 335436 234028 335442
rect 233976 335378 234028 335384
rect 233988 13326 234016 335378
rect 233976 13320 234028 13326
rect 233976 13262 234028 13268
rect 233884 12232 233936 12238
rect 233884 12174 233936 12180
rect 232504 11960 232556 11966
rect 232504 11902 232556 11908
rect 231032 8560 231084 8566
rect 231032 8502 231084 8508
rect 229836 7132 229888 7138
rect 229836 7074 229888 7080
rect 228732 4616 228784 4622
rect 228732 4558 228784 4564
rect 227628 4208 227680 4214
rect 227628 4150 227680 4156
rect 228744 480 228772 4558
rect 229848 480 229876 7074
rect 231044 480 231072 8502
rect 233424 7064 233476 7070
rect 233424 7006 233476 7012
rect 232228 4548 232280 4554
rect 232228 4490 232280 4496
rect 232240 480 232268 4490
rect 233436 480 233464 7006
rect 234632 6866 234660 457286
rect 240782 457328 240838 457337
rect 237250 457286 237360 457314
rect 238924 457298 239260 457314
rect 238924 457292 239272 457298
rect 238924 457286 239220 457292
rect 237194 457263 237250 457272
rect 240488 457286 240782 457314
rect 242346 457328 242402 457337
rect 242052 457286 242346 457314
rect 240782 457263 240838 457272
rect 243910 457328 243966 457337
rect 243616 457286 243910 457314
rect 242346 457263 242402 457272
rect 245474 457328 245530 457337
rect 245272 457286 245474 457314
rect 243910 457263 243966 457272
rect 246946 457328 247002 457337
rect 246836 457286 246946 457314
rect 245474 457263 245530 457272
rect 246946 457263 247002 457272
rect 248234 457328 248290 457337
rect 250258 457328 250314 457337
rect 248290 457286 248400 457314
rect 249964 457286 250258 457314
rect 248234 457263 248290 457272
rect 251822 457328 251878 457337
rect 251528 457286 251822 457314
rect 250258 457263 250314 457272
rect 253386 457328 253442 457337
rect 253092 457286 253386 457314
rect 251822 457263 251878 457272
rect 256514 457328 256570 457337
rect 254748 457298 255084 457314
rect 254748 457292 255096 457298
rect 254748 457286 255044 457292
rect 253386 457263 253442 457272
rect 239220 457234 239272 457240
rect 256312 457286 256514 457314
rect 256514 457263 256570 457272
rect 257526 457328 257582 457337
rect 259274 457328 259330 457337
rect 257582 457286 257876 457314
rect 257526 457263 257582 457272
rect 261298 457328 261354 457337
rect 259330 457286 259440 457314
rect 261004 457286 261298 457314
rect 259274 457263 259330 457272
rect 262862 457328 262918 457337
rect 262568 457286 262862 457314
rect 261298 457263 261354 457272
rect 264518 457328 264574 457337
rect 264224 457286 264518 457314
rect 262862 457263 262918 457272
rect 265788 457298 266124 457314
rect 275264 457298 275600 457314
rect 278392 457308 278688 457314
rect 278392 457302 278740 457308
rect 382278 457328 382334 457337
rect 265788 457292 266136 457298
rect 265788 457286 266084 457292
rect 264518 457263 264574 457272
rect 255044 457234 255096 457240
rect 275264 457292 275612 457298
rect 275264 457286 275560 457292
rect 266084 457234 266136 457240
rect 278392 457286 278728 457302
rect 384302 457328 384358 457337
rect 382334 457286 382628 457314
rect 384192 457286 384302 457314
rect 382278 457263 382334 457272
rect 384302 457263 384358 457272
rect 385406 457328 385462 457337
rect 387062 457328 387118 457337
rect 385462 457286 385756 457314
rect 385406 457263 385462 457272
rect 388626 457328 388682 457337
rect 387118 457286 387412 457314
rect 387062 457263 387118 457272
rect 390190 457328 390246 457337
rect 388682 457286 388976 457314
rect 388626 457263 388682 457272
rect 393502 457328 393558 457337
rect 390246 457286 390540 457314
rect 390190 457263 390246 457272
rect 394882 457328 394938 457337
rect 393558 457286 393668 457314
rect 393502 457263 393558 457272
rect 396538 457328 396594 457337
rect 394938 457286 395232 457314
rect 394882 457263 394938 457272
rect 398102 457328 398158 457337
rect 396594 457286 396888 457314
rect 396538 457263 396594 457272
rect 399666 457328 399722 457337
rect 398158 457286 398452 457314
rect 398102 457263 398158 457272
rect 401230 457328 401286 457337
rect 399722 457286 400016 457314
rect 399666 457263 399722 457272
rect 402978 457328 403034 457337
rect 401286 457286 401580 457314
rect 401230 457263 401286 457272
rect 404358 457328 404414 457337
rect 403034 457286 403144 457314
rect 402978 457263 403034 457272
rect 406014 457328 406070 457337
rect 404414 457286 404708 457314
rect 404358 457263 404414 457272
rect 409142 457328 409198 457337
rect 406070 457286 406364 457314
rect 406014 457263 406070 457272
rect 410706 457328 410762 457337
rect 409198 457286 409492 457314
rect 409142 457263 409198 457272
rect 412270 457328 412326 457337
rect 410762 457286 411056 457314
rect 410706 457263 410762 457272
rect 412326 457286 412620 457314
rect 414184 457286 414980 457314
rect 412270 457263 412326 457272
rect 275560 457234 275612 457240
rect 234724 338014 235152 338042
rect 235276 338014 235428 338042
rect 235552 338014 235796 338042
rect 234620 6860 234672 6866
rect 234620 6802 234672 6808
rect 234724 4826 234752 338014
rect 234804 330472 234856 330478
rect 234804 330414 234856 330420
rect 234816 4962 234844 330414
rect 235276 316034 235304 338014
rect 235552 330478 235580 338014
rect 236150 337770 236178 338028
rect 236288 338014 236532 338042
rect 236656 338014 236900 338042
rect 237024 338014 237268 338042
rect 237484 338014 237636 338042
rect 237760 338014 238004 338042
rect 238128 338014 238372 338042
rect 238496 338014 238740 338042
rect 238864 338014 239108 338042
rect 239232 338014 239476 338042
rect 239600 338014 239844 338042
rect 240152 338014 240212 338042
rect 240336 338014 240580 338042
rect 240704 338014 240948 338042
rect 241072 338014 241316 338042
rect 236150 337742 236224 337770
rect 235540 330472 235592 330478
rect 235540 330414 235592 330420
rect 236092 330472 236144 330478
rect 236092 330414 236144 330420
rect 234908 316006 235304 316034
rect 234804 4956 234856 4962
rect 234804 4898 234856 4904
rect 234908 4894 234936 316006
rect 234988 8492 235040 8498
rect 234988 8434 235040 8440
rect 234896 4888 234948 4894
rect 234896 4830 234948 4836
rect 234712 4820 234764 4826
rect 234712 4762 234764 4768
rect 235000 3482 235028 8434
rect 236104 5030 236132 330414
rect 236196 7614 236224 337742
rect 236288 336025 236316 338014
rect 236274 336016 236330 336025
rect 236274 335951 236330 335960
rect 236656 316034 236684 338014
rect 237024 330478 237052 338014
rect 237012 330472 237064 330478
rect 237012 330414 237064 330420
rect 237380 330472 237432 330478
rect 237380 330414 237432 330420
rect 236288 316006 236684 316034
rect 236184 7608 236236 7614
rect 236184 7550 236236 7556
rect 236092 5024 236144 5030
rect 236092 4966 236144 4972
rect 235816 4820 235868 4826
rect 235816 4762 235868 4768
rect 234632 3454 235028 3482
rect 234632 480 234660 3454
rect 235828 480 235856 4762
rect 236288 3369 236316 316006
rect 237392 7682 237420 330414
rect 237484 8974 237512 338014
rect 237760 327758 237788 338014
rect 238128 336161 238156 338014
rect 238114 336152 238170 336161
rect 238114 336087 238170 336096
rect 238496 330478 238524 338014
rect 238864 334626 238892 338014
rect 239232 335354 239260 338014
rect 238956 335326 239260 335354
rect 238852 334620 238904 334626
rect 238852 334562 238904 334568
rect 238956 330528 238984 335326
rect 238864 330500 238984 330528
rect 238484 330472 238536 330478
rect 238484 330414 238536 330420
rect 237748 327752 237800 327758
rect 237748 327694 237800 327700
rect 237472 8968 237524 8974
rect 237472 8910 237524 8916
rect 238116 8968 238168 8974
rect 238116 8910 238168 8916
rect 237380 7676 237432 7682
rect 237380 7618 237432 7624
rect 237012 7608 237064 7614
rect 237012 7550 237064 7556
rect 236274 3360 236330 3369
rect 236274 3295 236330 3304
rect 237024 480 237052 7550
rect 238128 480 238156 8910
rect 238864 3505 238892 330500
rect 239600 316034 239628 338014
rect 238956 316006 239628 316034
rect 238956 3641 238984 316006
rect 240152 7750 240180 338014
rect 240336 329118 240364 338014
rect 240704 336297 240732 338014
rect 241072 336433 241100 338014
rect 241670 337770 241698 338028
rect 241900 338014 242052 338042
rect 242176 338014 242420 338042
rect 242544 338014 242788 338042
rect 243004 338014 243156 338042
rect 243280 338014 243524 338042
rect 243648 338014 243892 338042
rect 244016 338014 244260 338042
rect 244476 338014 244628 338042
rect 244752 338014 244996 338042
rect 245120 338014 245364 338042
rect 245672 338014 245732 338042
rect 245856 338014 246100 338042
rect 246224 338014 246468 338042
rect 246592 338014 246836 338042
rect 247112 338014 247264 338042
rect 241670 337742 241744 337770
rect 241058 336424 241114 336433
rect 241058 336359 241114 336368
rect 240690 336288 240746 336297
rect 240690 336223 240746 336232
rect 241612 330540 241664 330546
rect 241612 330482 241664 330488
rect 240324 329112 240376 329118
rect 240324 329054 240376 329060
rect 240140 7744 240192 7750
rect 240140 7686 240192 7692
rect 240508 7676 240560 7682
rect 240508 7618 240560 7624
rect 239312 4888 239364 4894
rect 239312 4830 239364 4836
rect 238942 3632 238998 3641
rect 238942 3567 238998 3576
rect 238850 3496 238906 3505
rect 238850 3431 238906 3440
rect 239324 480 239352 4830
rect 240520 480 240548 7618
rect 241624 3466 241652 330482
rect 241716 8514 241744 337742
rect 241900 333266 241928 338014
rect 241888 333260 241940 333266
rect 241888 333202 241940 333208
rect 242176 316034 242204 338014
rect 242544 330546 242572 338014
rect 242532 330540 242584 330546
rect 242532 330482 242584 330488
rect 241808 316006 242204 316034
rect 241808 16574 241836 316006
rect 241808 16546 241928 16574
rect 241716 8486 241836 8514
rect 241704 8424 241756 8430
rect 241704 8366 241756 8372
rect 241612 3460 241664 3466
rect 241612 3402 241664 3408
rect 241716 480 241744 8366
rect 241808 7818 241836 8486
rect 241796 7812 241848 7818
rect 241796 7754 241848 7760
rect 241900 3777 241928 16546
rect 243004 7886 243032 338014
rect 243280 334694 243308 338014
rect 243648 336054 243676 338014
rect 243636 336048 243688 336054
rect 243636 335990 243688 335996
rect 243268 334688 243320 334694
rect 243268 334630 243320 334636
rect 244016 316034 244044 338014
rect 244476 331906 244504 338014
rect 244464 331900 244516 331906
rect 244464 331842 244516 331848
rect 244372 330540 244424 330546
rect 244372 330482 244424 330488
rect 243096 316006 244044 316034
rect 243096 7954 243124 316006
rect 244384 9042 244412 330482
rect 244752 316034 244780 338014
rect 245120 330546 245148 338014
rect 245108 330540 245160 330546
rect 245108 330482 245160 330488
rect 245672 330478 245700 338014
rect 245856 336122 245884 338014
rect 245844 336116 245896 336122
rect 245844 336058 245896 336064
rect 245660 330472 245712 330478
rect 245660 330414 245712 330420
rect 246224 316034 246252 338014
rect 246592 329186 246620 338014
rect 247132 330540 247184 330546
rect 247132 330482 247184 330488
rect 246580 329180 246632 329186
rect 246580 329122 246632 329128
rect 244476 316006 244780 316034
rect 245856 316006 246252 316034
rect 244372 9036 244424 9042
rect 244372 8978 244424 8984
rect 243084 7948 243136 7954
rect 243084 7890 243136 7896
rect 242992 7880 243044 7886
rect 242992 7822 243044 7828
rect 244096 7744 244148 7750
rect 244096 7686 244148 7692
rect 242900 4956 242952 4962
rect 242900 4898 242952 4904
rect 241886 3768 241942 3777
rect 241886 3703 241942 3712
rect 242912 480 242940 4898
rect 244108 480 244136 7686
rect 244476 3534 244504 316006
rect 245856 9110 245884 316006
rect 247144 10334 247172 330482
rect 247132 10328 247184 10334
rect 247132 10270 247184 10276
rect 245844 9104 245896 9110
rect 245844 9046 245896 9052
rect 245200 9036 245252 9042
rect 245200 8978 245252 8984
rect 244464 3528 244516 3534
rect 244464 3470 244516 3476
rect 245212 480 245240 8978
rect 246396 5024 246448 5030
rect 246396 4966 246448 4972
rect 246408 480 246436 4966
rect 247236 3602 247264 338014
rect 247328 338014 247480 338042
rect 247604 338014 247848 338042
rect 247972 338014 248216 338042
rect 247328 330546 247356 338014
rect 247604 333334 247632 338014
rect 247972 336190 248000 338014
rect 248570 337770 248598 338028
rect 248708 338014 248952 338042
rect 249076 338014 249320 338042
rect 249444 338014 249688 338042
rect 249996 338014 250056 338042
rect 250180 338014 250424 338042
rect 250548 338014 250792 338042
rect 250916 338014 251160 338042
rect 251284 338014 251528 338042
rect 251652 338014 251896 338042
rect 252020 338014 252264 338042
rect 252572 338014 252632 338042
rect 252756 338014 253000 338042
rect 253124 338014 253368 338042
rect 253492 338014 253736 338042
rect 248570 337742 248644 337770
rect 247960 336184 248012 336190
rect 247960 336126 248012 336132
rect 247592 333328 247644 333334
rect 247592 333270 247644 333276
rect 247316 330540 247368 330546
rect 247316 330482 247368 330488
rect 248512 330540 248564 330546
rect 248512 330482 248564 330488
rect 247592 7812 247644 7818
rect 247592 7754 247644 7760
rect 247224 3596 247276 3602
rect 247224 3538 247276 3544
rect 247604 480 247632 7754
rect 248524 6186 248552 330482
rect 248616 10402 248644 337742
rect 248708 330614 248736 338014
rect 248696 330608 248748 330614
rect 248696 330550 248748 330556
rect 249076 316034 249104 338014
rect 249444 330546 249472 338014
rect 249432 330540 249484 330546
rect 249432 330482 249484 330488
rect 249892 330540 249944 330546
rect 249892 330482 249944 330488
rect 248708 316006 249104 316034
rect 248604 10396 248656 10402
rect 248604 10338 248656 10344
rect 248512 6180 248564 6186
rect 248512 6122 248564 6128
rect 248708 3670 248736 316006
rect 249904 10538 249932 330482
rect 249892 10532 249944 10538
rect 249892 10474 249944 10480
rect 249996 10470 250024 338014
rect 250180 331974 250208 338014
rect 250168 331968 250220 331974
rect 250168 331910 250220 331916
rect 250548 316034 250576 338014
rect 250916 330546 250944 338014
rect 251284 336258 251312 338014
rect 251272 336252 251324 336258
rect 251272 336194 251324 336200
rect 250904 330540 250956 330546
rect 250904 330482 250956 330488
rect 251272 330540 251324 330546
rect 251272 330482 251324 330488
rect 250088 316006 250576 316034
rect 249984 10464 250036 10470
rect 249984 10406 250036 10412
rect 248788 9104 248840 9110
rect 248788 9046 248840 9052
rect 248696 3664 248748 3670
rect 248696 3606 248748 3612
rect 248800 480 248828 9046
rect 250088 6254 250116 316006
rect 251088 11960 251140 11966
rect 251088 11902 251140 11908
rect 250076 6248 250128 6254
rect 250076 6190 250128 6196
rect 251100 3534 251128 11902
rect 251284 10606 251312 330482
rect 251652 316034 251680 338014
rect 252020 330546 252048 338014
rect 252008 330540 252060 330546
rect 252008 330482 252060 330488
rect 252572 329254 252600 338014
rect 252756 336682 252784 338014
rect 252664 336654 252784 336682
rect 252560 329248 252612 329254
rect 252560 329190 252612 329196
rect 251376 316006 251680 316034
rect 251272 10600 251324 10606
rect 251272 10542 251324 10548
rect 251180 7948 251232 7954
rect 251180 7890 251232 7896
rect 249984 3528 250036 3534
rect 249984 3470 250036 3476
rect 251088 3528 251140 3534
rect 251088 3470 251140 3476
rect 249996 480 250024 3470
rect 251192 480 251220 7890
rect 251376 6322 251404 316006
rect 252376 14476 252428 14482
rect 252376 14418 252428 14424
rect 251364 6316 251416 6322
rect 251364 6258 251416 6264
rect 252388 480 252416 14418
rect 252664 6390 252692 336654
rect 253124 335354 253152 338014
rect 252756 335326 253152 335354
rect 252756 10674 252784 335326
rect 253492 316034 253520 338014
rect 254090 337770 254118 338028
rect 254228 338014 254472 338042
rect 254596 338014 254840 338042
rect 254964 338014 255208 338042
rect 255516 338014 255576 338042
rect 255700 338014 255944 338042
rect 256068 338014 256312 338042
rect 256436 338014 256680 338042
rect 256804 338014 257048 338042
rect 257172 338014 257416 338042
rect 257540 338014 257784 338042
rect 258092 338014 258152 338042
rect 258276 338014 258520 338042
rect 258644 338014 258888 338042
rect 259012 338014 259164 338042
rect 254090 337742 254164 337770
rect 253940 330540 253992 330546
rect 253940 330482 253992 330488
rect 252848 316006 253520 316034
rect 252744 10668 252796 10674
rect 252744 10610 252796 10616
rect 252652 6384 252704 6390
rect 252652 6326 252704 6332
rect 252848 3738 252876 316006
rect 253480 10600 253532 10606
rect 253480 10542 253532 10548
rect 252836 3732 252888 3738
rect 252836 3674 252888 3680
rect 253492 480 253520 10542
rect 253952 3806 253980 330482
rect 254032 330472 254084 330478
rect 254032 330414 254084 330420
rect 254044 6526 254072 330414
rect 254032 6520 254084 6526
rect 254032 6462 254084 6468
rect 254136 6458 254164 337742
rect 254228 10742 254256 338014
rect 254596 330546 254624 338014
rect 254584 330540 254636 330546
rect 254584 330482 254636 330488
rect 254964 330478 254992 338014
rect 255412 330540 255464 330546
rect 255412 330482 255464 330488
rect 254952 330472 255004 330478
rect 254952 330414 255004 330420
rect 255320 329656 255372 329662
rect 255320 329598 255372 329604
rect 254216 10736 254268 10742
rect 254216 10678 254268 10684
rect 254676 7880 254728 7886
rect 254676 7822 254728 7828
rect 254124 6452 254176 6458
rect 254124 6394 254176 6400
rect 253940 3800 253992 3806
rect 253940 3742 253992 3748
rect 254688 480 254716 7822
rect 255332 3874 255360 329598
rect 255424 6594 255452 330482
rect 255516 10810 255544 338014
rect 255700 329662 255728 338014
rect 256068 330546 256096 338014
rect 256056 330540 256108 330546
rect 256056 330482 256108 330488
rect 255688 329656 255740 329662
rect 255688 329598 255740 329604
rect 256436 316034 256464 338014
rect 256804 336682 256832 338014
rect 255608 316006 256464 316034
rect 256712 336654 256832 336682
rect 255608 10878 255636 316006
rect 255596 10872 255648 10878
rect 255596 10814 255648 10820
rect 255504 10804 255556 10810
rect 255504 10746 255556 10752
rect 256608 10328 256660 10334
rect 256608 10270 256660 10276
rect 255412 6588 255464 6594
rect 255412 6530 255464 6536
rect 255320 3868 255372 3874
rect 255320 3810 255372 3816
rect 256620 3534 256648 10270
rect 256712 3942 256740 336654
rect 257172 335354 257200 338014
rect 256804 335326 257200 335354
rect 256804 8022 256832 335326
rect 257540 316034 257568 338014
rect 256896 316006 257568 316034
rect 256896 11762 256924 316006
rect 256884 11756 256936 11762
rect 256884 11698 256936 11704
rect 256792 8016 256844 8022
rect 256792 7958 256844 7964
rect 257068 6180 257120 6186
rect 257068 6122 257120 6128
rect 256700 3936 256752 3942
rect 256700 3878 256752 3884
rect 255872 3528 255924 3534
rect 255872 3470 255924 3476
rect 256608 3528 256660 3534
rect 256608 3470 256660 3476
rect 255884 480 255912 3470
rect 257080 480 257108 6122
rect 258092 4010 258120 338014
rect 258172 330540 258224 330546
rect 258172 330482 258224 330488
rect 258184 4078 258212 330482
rect 258276 8242 258304 338014
rect 258644 316034 258672 338014
rect 259012 330546 259040 338014
rect 259518 337770 259546 338028
rect 259656 338014 259900 338042
rect 260024 338014 260268 338042
rect 260392 338014 260636 338042
rect 260944 338014 261004 338042
rect 261128 338014 261372 338042
rect 261496 338014 261740 338042
rect 261956 338014 262108 338042
rect 259518 337742 259592 337770
rect 259460 336252 259512 336258
rect 259460 336194 259512 336200
rect 259472 334762 259500 336194
rect 259460 334756 259512 334762
rect 259460 334698 259512 334704
rect 259000 330540 259052 330546
rect 259000 330482 259052 330488
rect 258368 316006 258672 316034
rect 258368 11830 258396 316006
rect 258356 11824 258408 11830
rect 258356 11766 258408 11772
rect 258276 8214 258396 8242
rect 258368 8158 258396 8214
rect 259564 8158 259592 337742
rect 259656 330682 259684 338014
rect 259644 330676 259696 330682
rect 259644 330618 259696 330624
rect 260024 316034 260052 338014
rect 260392 333402 260420 338014
rect 260944 334830 260972 338014
rect 260932 334824 260984 334830
rect 260932 334766 260984 334772
rect 260380 333396 260432 333402
rect 260380 333338 260432 333344
rect 261128 316034 261156 338014
rect 261496 336258 261524 338014
rect 261484 336252 261536 336258
rect 261484 336194 261536 336200
rect 261956 333470 261984 338014
rect 262462 337770 262490 338028
rect 262600 338014 262844 338042
rect 262968 338014 263212 338042
rect 263336 338014 263580 338042
rect 263704 338014 263948 338042
rect 264072 338014 264316 338042
rect 264440 338014 264684 338042
rect 262462 337742 262536 337770
rect 261944 333464 261996 333470
rect 261944 333406 261996 333412
rect 262404 330540 262456 330546
rect 262404 330482 262456 330488
rect 262312 330472 262364 330478
rect 262312 330414 262364 330420
rect 259748 316006 260052 316034
rect 261036 316006 261156 316034
rect 258356 8152 258408 8158
rect 258356 8094 258408 8100
rect 259552 8152 259604 8158
rect 259552 8094 259604 8100
rect 258264 8084 258316 8090
rect 258264 8026 258316 8032
rect 258172 4072 258224 4078
rect 258172 4014 258224 4020
rect 258080 4004 258132 4010
rect 258080 3946 258132 3952
rect 258276 480 258304 8026
rect 259460 6316 259512 6322
rect 259460 6258 259512 6264
rect 259472 480 259500 6258
rect 259748 4146 259776 316006
rect 260656 10668 260708 10674
rect 260656 10610 260708 10616
rect 259736 4140 259788 4146
rect 259736 4082 259788 4088
rect 260668 480 260696 10610
rect 261036 3398 261064 316006
rect 261760 8084 261812 8090
rect 261760 8026 261812 8032
rect 261024 3392 261076 3398
rect 261024 3334 261076 3340
rect 261772 480 261800 8026
rect 262324 3262 262352 330414
rect 262416 10946 262444 330482
rect 262404 10940 262456 10946
rect 262404 10882 262456 10888
rect 262508 3330 262536 337742
rect 262600 330546 262628 338014
rect 262968 333538 262996 338014
rect 262956 333532 263008 333538
rect 262956 333474 263008 333480
rect 262588 330540 262640 330546
rect 262588 330482 262640 330488
rect 263336 330478 263364 338014
rect 263508 336048 263560 336054
rect 263508 335990 263560 335996
rect 263324 330472 263376 330478
rect 263324 330414 263376 330420
rect 263520 3534 263548 335990
rect 263704 11014 263732 338014
rect 264072 332042 264100 338014
rect 264060 332036 264112 332042
rect 264060 331978 264112 331984
rect 264440 316034 264468 338014
rect 265038 337770 265066 338028
rect 265176 338014 265420 338042
rect 265544 338014 265788 338042
rect 265912 338014 266156 338042
rect 266372 338014 266524 338042
rect 266648 338014 266892 338042
rect 267016 338014 267260 338042
rect 267384 338014 267628 338042
rect 267844 338014 267996 338042
rect 268120 338014 268364 338042
rect 268488 338014 268732 338042
rect 268856 338014 269100 338042
rect 269316 338014 269468 338042
rect 269592 338014 269836 338042
rect 269960 338014 270204 338042
rect 270572 338014 270724 338042
rect 265038 337742 265112 337770
rect 264520 336252 264572 336258
rect 264520 336194 264572 336200
rect 264532 332110 264560 336194
rect 264520 332104 264572 332110
rect 264520 332046 264572 332052
rect 263796 316006 264468 316034
rect 263692 11008 263744 11014
rect 263692 10950 263744 10956
rect 262956 3528 263008 3534
rect 262956 3470 263008 3476
rect 263508 3528 263560 3534
rect 263508 3470 263560 3476
rect 262496 3324 262548 3330
rect 262496 3266 262548 3272
rect 262312 3256 262364 3262
rect 262312 3198 262364 3204
rect 262968 480 262996 3470
rect 263796 3194 263824 316006
rect 264888 10396 264940 10402
rect 264888 10338 264940 10344
rect 264900 3534 264928 10338
rect 265084 10266 265112 337742
rect 265176 336258 265204 338014
rect 265164 336252 265216 336258
rect 265164 336194 265216 336200
rect 265164 330540 265216 330546
rect 265164 330482 265216 330488
rect 265072 10260 265124 10266
rect 265072 10202 265124 10208
rect 265176 10198 265204 330482
rect 265544 316034 265572 338014
rect 265912 330546 265940 338014
rect 266372 332178 266400 338014
rect 266360 332172 266412 332178
rect 266360 332114 266412 332120
rect 265900 330540 265952 330546
rect 265900 330482 265952 330488
rect 266452 330540 266504 330546
rect 266452 330482 266504 330488
rect 265268 316006 265572 316034
rect 265164 10192 265216 10198
rect 265164 10134 265216 10140
rect 264152 3528 264204 3534
rect 264152 3470 264204 3476
rect 264888 3528 264940 3534
rect 264888 3470 264940 3476
rect 263784 3188 263836 3194
rect 263784 3130 263836 3136
rect 264164 480 264192 3470
rect 265268 3126 265296 316006
rect 266464 10130 266492 330482
rect 266452 10124 266504 10130
rect 266452 10066 266504 10072
rect 265348 8152 265400 8158
rect 265348 8094 265400 8100
rect 265256 3120 265308 3126
rect 265256 3062 265308 3068
rect 265360 480 265388 8094
rect 266544 3528 266596 3534
rect 266544 3470 266596 3476
rect 266556 480 266584 3470
rect 266648 3058 266676 338014
rect 267016 330546 267044 338014
rect 267384 330750 267412 338014
rect 267844 336326 267872 338014
rect 267832 336320 267884 336326
rect 267832 336262 267884 336268
rect 267648 336184 267700 336190
rect 267648 336126 267700 336132
rect 267372 330744 267424 330750
rect 267372 330686 267424 330692
rect 267004 330540 267056 330546
rect 267004 330482 267056 330488
rect 267660 3534 267688 336126
rect 267740 335368 267792 335374
rect 268120 335354 268148 338014
rect 267740 335310 267792 335316
rect 267936 335326 268148 335354
rect 267752 329458 267780 335310
rect 267936 330562 267964 335326
rect 268488 330818 268516 338014
rect 268476 330812 268528 330818
rect 268476 330754 268528 330760
rect 267844 330534 267964 330562
rect 267740 329452 267792 329458
rect 267740 329394 267792 329400
rect 267844 10062 267872 330534
rect 268856 316034 268884 338014
rect 267936 316006 268884 316034
rect 267832 10056 267884 10062
rect 267832 9998 267884 10004
rect 267648 3528 267700 3534
rect 267648 3470 267700 3476
rect 267740 3460 267792 3466
rect 267740 3402 267792 3408
rect 266636 3052 266688 3058
rect 266636 2994 266688 3000
rect 267752 480 267780 3402
rect 267936 2990 267964 316006
rect 269028 10464 269080 10470
rect 269028 10406 269080 10412
rect 268844 6248 268896 6254
rect 268844 6190 268896 6196
rect 267924 2984 267976 2990
rect 267924 2926 267976 2932
rect 268856 480 268884 6190
rect 269040 3466 269068 10406
rect 269316 9994 269344 338014
rect 269592 329322 269620 338014
rect 269960 336394 269988 338014
rect 269948 336388 270000 336394
rect 269948 336330 270000 336336
rect 270040 336252 270092 336258
rect 270040 336194 270092 336200
rect 270052 329390 270080 336194
rect 270408 336116 270460 336122
rect 270408 336058 270460 336064
rect 270040 329384 270092 329390
rect 270040 329326 270092 329332
rect 269580 329316 269632 329322
rect 269580 329258 269632 329264
rect 269304 9988 269356 9994
rect 269304 9930 269356 9936
rect 270420 6914 270448 336058
rect 270592 330540 270644 330546
rect 270592 330482 270644 330488
rect 270604 9858 270632 330482
rect 270696 9926 270724 338014
rect 270880 338014 270940 338042
rect 271064 338014 271216 338042
rect 271340 338014 271584 338042
rect 271892 338014 271952 338042
rect 272076 338014 272320 338042
rect 272444 338014 272688 338042
rect 272812 338014 273056 338042
rect 273272 338014 273424 338042
rect 273548 338014 273792 338042
rect 273916 338014 274160 338042
rect 274284 338014 274528 338042
rect 274744 338014 274896 338042
rect 275020 338014 275264 338042
rect 275388 338014 275632 338042
rect 275756 338014 276000 338042
rect 276216 338014 276368 338042
rect 276492 338014 276736 338042
rect 276860 338014 277104 338042
rect 270880 330886 270908 338014
rect 270868 330880 270920 330886
rect 270868 330822 270920 330828
rect 271064 316034 271092 338014
rect 271340 330546 271368 338014
rect 271892 336258 271920 338014
rect 271880 336252 271932 336258
rect 271880 336194 271932 336200
rect 271328 330540 271380 330546
rect 271328 330482 271380 330488
rect 271972 329860 272024 329866
rect 271972 329802 272024 329808
rect 270788 316006 271092 316034
rect 270684 9920 270736 9926
rect 270684 9862 270736 9868
rect 270592 9852 270644 9858
rect 270592 9794 270644 9800
rect 270052 6886 270448 6914
rect 269028 3460 269080 3466
rect 269028 3402 269080 3408
rect 270052 480 270080 6886
rect 270788 2922 270816 316006
rect 271788 10532 271840 10538
rect 271788 10474 271840 10480
rect 271800 3534 271828 10474
rect 271984 9790 272012 329802
rect 271972 9784 272024 9790
rect 271972 9726 272024 9732
rect 271236 3528 271288 3534
rect 271236 3470 271288 3476
rect 271788 3528 271840 3534
rect 271788 3470 271840 3476
rect 270776 2916 270828 2922
rect 270776 2858 270828 2864
rect 271248 480 271276 3470
rect 272076 2854 272104 338014
rect 272444 329866 272472 338014
rect 272812 335374 272840 338014
rect 273272 336462 273300 338014
rect 273260 336456 273312 336462
rect 273260 336398 273312 336404
rect 273548 335442 273576 338014
rect 273916 335646 273944 338014
rect 273904 335640 273956 335646
rect 273904 335582 273956 335588
rect 273536 335436 273588 335442
rect 273536 335378 273588 335384
rect 272800 335368 272852 335374
rect 272800 335310 272852 335316
rect 272432 329860 272484 329866
rect 272432 329802 272484 329808
rect 274284 316034 274312 338014
rect 274548 336252 274600 336258
rect 274548 336194 274600 336200
rect 274456 335368 274508 335374
rect 274456 335310 274508 335316
rect 274468 332246 274496 335310
rect 274456 332240 274508 332246
rect 274456 332182 274508 332188
rect 273456 316006 274312 316034
rect 273456 13122 273484 316006
rect 273444 13116 273496 13122
rect 273444 13058 273496 13064
rect 274560 3534 274588 336194
rect 274640 326392 274692 326398
rect 274640 326334 274692 326340
rect 274652 5166 274680 326334
rect 274640 5160 274692 5166
rect 274640 5102 274692 5108
rect 274744 5098 274772 338014
rect 275020 335354 275048 338014
rect 274836 335326 275048 335354
rect 274836 6662 274864 335326
rect 275388 316034 275416 338014
rect 275756 326398 275784 338014
rect 276020 336456 276072 336462
rect 276020 336398 276072 336404
rect 276032 335034 276060 336398
rect 276020 335028 276072 335034
rect 276020 334970 276072 334976
rect 276216 326466 276244 338014
rect 276492 335354 276520 338014
rect 276860 335986 276888 338014
rect 277458 337770 277486 338028
rect 277596 338014 277840 338042
rect 277964 338014 278208 338042
rect 278332 338014 278576 338042
rect 278792 338014 278944 338042
rect 279068 338014 279312 338042
rect 279436 338014 279680 338042
rect 279804 338014 280048 338042
rect 280264 338014 280416 338042
rect 280540 338014 280784 338042
rect 280908 338014 281152 338042
rect 281460 338014 281520 338042
rect 281736 338014 281888 338042
rect 282012 338014 282256 338042
rect 282380 338014 282624 338042
rect 277458 337742 277532 337770
rect 277308 336388 277360 336394
rect 277308 336330 277360 336336
rect 276848 335980 276900 335986
rect 276848 335922 276900 335928
rect 276308 335326 276520 335354
rect 276204 326460 276256 326466
rect 276204 326402 276256 326408
rect 275744 326392 275796 326398
rect 275744 326334 275796 326340
rect 276204 326256 276256 326262
rect 276204 326198 276256 326204
rect 276112 323672 276164 323678
rect 276112 323614 276164 323620
rect 274928 316006 275416 316034
rect 274928 9178 274956 316006
rect 276124 9246 276152 323614
rect 276112 9240 276164 9246
rect 276112 9182 276164 9188
rect 274916 9172 274968 9178
rect 274916 9114 274968 9120
rect 276216 8226 276244 326198
rect 276308 323678 276336 335326
rect 276296 323672 276348 323678
rect 276296 323614 276348 323620
rect 276204 8220 276256 8226
rect 276204 8162 276256 8168
rect 274824 6656 274876 6662
rect 274824 6598 274876 6604
rect 274732 5092 274784 5098
rect 274732 5034 274784 5040
rect 274824 5092 274876 5098
rect 274824 5034 274876 5040
rect 273628 3528 273680 3534
rect 273628 3470 273680 3476
rect 274548 3528 274600 3534
rect 274548 3470 274600 3476
rect 272432 3460 272484 3466
rect 272432 3402 272484 3408
rect 272064 2848 272116 2854
rect 272064 2790 272116 2796
rect 272444 480 272472 3402
rect 273640 480 273668 3470
rect 274836 480 274864 5034
rect 277320 3534 277348 336330
rect 277400 336320 277452 336326
rect 277400 336262 277452 336268
rect 277412 330954 277440 336262
rect 277400 330948 277452 330954
rect 277400 330890 277452 330896
rect 277504 326398 277532 337742
rect 277492 326392 277544 326398
rect 277492 326334 277544 326340
rect 277492 325168 277544 325174
rect 277492 325110 277544 325116
rect 277504 7546 277532 325110
rect 277596 15910 277624 338014
rect 277964 334898 277992 338014
rect 277952 334892 278004 334898
rect 277952 334834 278004 334840
rect 277676 326392 277728 326398
rect 277676 326334 277728 326340
rect 277584 15904 277636 15910
rect 277584 15846 277636 15852
rect 277688 8294 277716 326334
rect 278332 325174 278360 338014
rect 278792 335374 278820 338014
rect 279068 336462 279096 338014
rect 279056 336456 279108 336462
rect 279056 336398 279108 336404
rect 278780 335368 278832 335374
rect 278780 335310 278832 335316
rect 278320 325168 278372 325174
rect 278320 325110 278372 325116
rect 279436 316034 279464 338014
rect 279804 336326 279832 338014
rect 279792 336320 279844 336326
rect 279792 336262 279844 336268
rect 280264 334966 280292 338014
rect 280252 334960 280304 334966
rect 280252 334902 280304 334908
rect 280252 326392 280304 326398
rect 280252 326334 280304 326340
rect 278976 316006 279464 316034
rect 277676 8288 277728 8294
rect 277676 8230 277728 8236
rect 277492 7540 277544 7546
rect 277492 7482 277544 7488
rect 278976 7478 279004 316006
rect 280264 13190 280292 326334
rect 280540 316034 280568 338014
rect 280908 326398 280936 338014
rect 281356 335980 281408 335986
rect 281356 335922 281408 335928
rect 281368 331214 281396 335922
rect 281460 333606 281488 338014
rect 281448 333600 281500 333606
rect 281448 333542 281500 333548
rect 281368 331186 281488 331214
rect 280896 326392 280948 326398
rect 280896 326334 280948 326340
rect 280356 316006 280568 316034
rect 280252 13184 280304 13190
rect 280252 13126 280304 13132
rect 278964 7472 279016 7478
rect 278964 7414 279016 7420
rect 280356 7410 280384 316006
rect 280344 7404 280396 7410
rect 280344 7346 280396 7352
rect 278320 5160 278372 5166
rect 278320 5102 278372 5108
rect 276020 3528 276072 3534
rect 276020 3470 276072 3476
rect 277308 3528 277360 3534
rect 277308 3470 277360 3476
rect 276032 480 276060 3470
rect 277122 3360 277178 3369
rect 277122 3295 277178 3304
rect 277136 480 277164 3295
rect 278332 480 278360 5102
rect 279516 3596 279568 3602
rect 279516 3538 279568 3544
rect 279528 480 279556 3538
rect 281460 3534 281488 331186
rect 281736 7342 281764 338014
rect 282012 331022 282040 338014
rect 282184 336320 282236 336326
rect 282184 336262 282236 336268
rect 282000 331016 282052 331022
rect 282000 330958 282052 330964
rect 282196 18630 282224 336262
rect 282380 335510 282408 338014
rect 282978 337770 283006 338028
rect 283116 338014 283268 338042
rect 283392 338014 283636 338042
rect 283760 338014 284004 338042
rect 282978 337742 283052 337770
rect 282644 336456 282696 336462
rect 282644 336398 282696 336404
rect 282368 335504 282420 335510
rect 282368 335446 282420 335452
rect 282656 333674 282684 336398
rect 282644 333668 282696 333674
rect 282644 333610 282696 333616
rect 282184 18624 282236 18630
rect 282184 18566 282236 18572
rect 281724 7336 281776 7342
rect 281724 7278 281776 7284
rect 283024 7274 283052 337742
rect 283116 336326 283144 338014
rect 283392 336462 283420 338014
rect 283380 336456 283432 336462
rect 283380 336398 283432 336404
rect 283104 336320 283156 336326
rect 283104 336262 283156 336268
rect 283760 316034 283788 338014
rect 284358 337770 284386 338028
rect 284496 338014 284740 338042
rect 284864 338014 285108 338042
rect 285232 338014 285476 338042
rect 285692 338014 285844 338042
rect 285968 338014 286212 338042
rect 286336 338014 286580 338042
rect 286704 338014 286948 338042
rect 287256 338014 287316 338042
rect 287440 338014 287684 338042
rect 287808 338014 288052 338042
rect 288176 338014 288420 338042
rect 288636 338014 288788 338042
rect 288912 338014 289156 338042
rect 289280 338014 289524 338042
rect 289832 338014 289892 338042
rect 290016 338014 290260 338042
rect 290384 338014 290628 338042
rect 290844 338014 290996 338042
rect 291212 338014 291364 338042
rect 291488 338014 291732 338042
rect 291856 338014 292100 338042
rect 292224 338014 292468 338042
rect 292684 338014 292836 338042
rect 292960 338014 293204 338042
rect 293328 338014 293572 338042
rect 293696 338014 293940 338042
rect 294156 338014 294308 338042
rect 294432 338014 294676 338042
rect 294800 338014 295044 338042
rect 295168 338014 295320 338042
rect 295444 338014 295688 338042
rect 295812 338014 296056 338042
rect 296180 338014 296424 338042
rect 296732 338014 296792 338042
rect 296916 338014 297160 338042
rect 297284 338014 297528 338042
rect 297652 338014 297896 338042
rect 298112 338014 298264 338042
rect 298388 338014 298632 338042
rect 298756 338014 299000 338042
rect 299124 338014 299368 338042
rect 299676 338014 299736 338042
rect 299860 338014 300104 338042
rect 300228 338014 300472 338042
rect 300596 338014 300840 338042
rect 301056 338014 301208 338042
rect 301332 338014 301576 338042
rect 301700 338014 301944 338042
rect 284358 337742 284432 337770
rect 283116 316006 283788 316034
rect 283012 7268 283064 7274
rect 283012 7210 283064 7216
rect 283116 7206 283144 316006
rect 284404 17270 284432 337742
rect 284496 335102 284524 338014
rect 284484 335096 284536 335102
rect 284484 335038 284536 335044
rect 284864 333742 284892 338014
rect 284852 333736 284904 333742
rect 284852 333678 284904 333684
rect 285232 316034 285260 338014
rect 285692 335578 285720 338014
rect 285680 335572 285732 335578
rect 285680 335514 285732 335520
rect 285772 330540 285824 330546
rect 285772 330482 285824 330488
rect 284496 316006 285260 316034
rect 284392 17264 284444 17270
rect 284392 17206 284444 17212
rect 284496 13258 284524 316006
rect 284484 13252 284536 13258
rect 284484 13194 284536 13200
rect 285784 11898 285812 330482
rect 285968 316034 285996 338014
rect 286336 330546 286364 338014
rect 286416 335980 286468 335986
rect 286416 335922 286468 335928
rect 286324 330540 286376 330546
rect 286324 330482 286376 330488
rect 286428 316034 286456 335922
rect 286704 335170 286732 338014
rect 286692 335164 286744 335170
rect 286692 335106 286744 335112
rect 287152 330540 287204 330546
rect 287152 330482 287204 330488
rect 285876 316006 285996 316034
rect 286336 316006 286456 316034
rect 285772 11892 285824 11898
rect 285772 11834 285824 11840
rect 283104 7200 283156 7206
rect 283104 7142 283156 7148
rect 285876 6730 285904 316006
rect 286336 10674 286364 316006
rect 286324 10668 286376 10674
rect 286324 10610 286376 10616
rect 285864 6724 285916 6730
rect 285864 6666 285916 6672
rect 287164 6118 287192 330482
rect 287256 6798 287284 338014
rect 287440 332314 287468 338014
rect 287808 335782 287836 338014
rect 287796 335776 287848 335782
rect 287796 335718 287848 335724
rect 287428 332308 287480 332314
rect 287428 332250 287480 332256
rect 288176 330546 288204 338014
rect 288532 336728 288584 336734
rect 288532 336670 288584 336676
rect 288440 336660 288492 336666
rect 288440 336602 288492 336608
rect 288348 335640 288400 335646
rect 288348 335582 288400 335588
rect 288164 330540 288216 330546
rect 288164 330482 288216 330488
rect 287244 6792 287296 6798
rect 287244 6734 287296 6740
rect 287152 6112 287204 6118
rect 287152 6054 287204 6060
rect 281908 4480 281960 4486
rect 281908 4422 281960 4428
rect 280712 3528 280764 3534
rect 280712 3470 280764 3476
rect 281448 3528 281500 3534
rect 281448 3470 281500 3476
rect 280724 480 280752 3470
rect 281920 480 281948 4422
rect 285404 4412 285456 4418
rect 285404 4354 285456 4360
rect 284300 3664 284352 3670
rect 284300 3606 284352 3612
rect 283102 3496 283158 3505
rect 283102 3431 283158 3440
rect 283116 480 283144 3431
rect 284312 480 284340 3606
rect 285416 480 285444 4354
rect 286600 3596 286652 3602
rect 286600 3538 286652 3544
rect 286612 480 286640 3538
rect 288360 3398 288388 335582
rect 288452 335238 288480 336602
rect 288440 335232 288492 335238
rect 288440 335174 288492 335180
rect 288544 333810 288572 336670
rect 288532 333804 288584 333810
rect 288532 333746 288584 333752
rect 288636 332382 288664 338014
rect 288912 335714 288940 338014
rect 289280 336682 289308 338014
rect 289832 336734 289860 338014
rect 289004 336654 289308 336682
rect 289820 336728 289872 336734
rect 289820 336670 289872 336676
rect 290016 336666 290044 338014
rect 290004 336660 290056 336666
rect 288900 335708 288952 335714
rect 288900 335650 288952 335656
rect 288624 332376 288676 332382
rect 288624 332318 288676 332324
rect 289004 316034 289032 336654
rect 290004 336602 290056 336608
rect 289084 335776 289136 335782
rect 289084 335718 289136 335724
rect 288636 316006 289032 316034
rect 288636 6050 288664 316006
rect 289096 10606 289124 335718
rect 290384 316034 290412 338014
rect 290844 332450 290872 338014
rect 291212 335918 291240 338014
rect 291384 336728 291436 336734
rect 291384 336670 291436 336676
rect 291200 335912 291252 335918
rect 291200 335854 291252 335860
rect 291396 332518 291424 336670
rect 291384 332512 291436 332518
rect 291384 332454 291436 332460
rect 290832 332444 290884 332450
rect 290832 332386 290884 332392
rect 291292 330540 291344 330546
rect 291292 330482 291344 330488
rect 290016 316006 290412 316034
rect 289084 10600 289136 10606
rect 289084 10542 289136 10548
rect 288624 6044 288676 6050
rect 288624 5986 288676 5992
rect 290016 5982 290044 316006
rect 291304 13394 291332 330482
rect 291488 316034 291516 338014
rect 291856 330546 291884 338014
rect 292224 336598 292252 338014
rect 292212 336592 292264 336598
rect 292212 336534 292264 336540
rect 291936 335912 291988 335918
rect 291936 335854 291988 335860
rect 291844 330540 291896 330546
rect 291844 330482 291896 330488
rect 291948 316034 291976 335854
rect 291396 316006 291516 316034
rect 291856 316006 291976 316034
rect 291292 13388 291344 13394
rect 291292 13330 291344 13336
rect 290004 5976 290056 5982
rect 290004 5918 290056 5924
rect 291396 5914 291424 316006
rect 291856 11966 291884 316006
rect 291844 11960 291896 11966
rect 291844 11902 291896 11908
rect 291384 5908 291436 5914
rect 291384 5850 291436 5856
rect 292684 5846 292712 338014
rect 292960 336734 292988 338014
rect 292948 336728 293000 336734
rect 292948 336670 293000 336676
rect 293328 336462 293356 338014
rect 293316 336456 293368 336462
rect 293316 336398 293368 336404
rect 293696 316034 293724 338014
rect 294052 330540 294104 330546
rect 294052 330482 294104 330488
rect 292776 316006 293724 316034
rect 292672 5840 292724 5846
rect 292672 5782 292724 5788
rect 292776 5778 292804 316006
rect 294064 9382 294092 330482
rect 294052 9376 294104 9382
rect 294052 9318 294104 9324
rect 294156 9314 294184 338014
rect 294432 336666 294460 338014
rect 294420 336660 294472 336666
rect 294420 336602 294472 336608
rect 294800 316034 294828 338014
rect 295168 330546 295196 338014
rect 295444 335374 295472 338014
rect 295432 335368 295484 335374
rect 295432 335310 295484 335316
rect 295812 333878 295840 338014
rect 296180 336682 296208 338014
rect 295904 336654 296208 336682
rect 296536 336660 296588 336666
rect 295800 333872 295852 333878
rect 295800 333814 295852 333820
rect 295156 330540 295208 330546
rect 295156 330482 295208 330488
rect 295904 316034 295932 336654
rect 296536 336602 296588 336608
rect 295984 335708 296036 335714
rect 295984 335650 296036 335656
rect 294248 316006 294828 316034
rect 295536 316006 295932 316034
rect 294144 9308 294196 9314
rect 294144 9250 294196 9256
rect 292764 5772 292816 5778
rect 292764 5714 292816 5720
rect 294248 5710 294276 316006
rect 295536 9450 295564 316006
rect 295524 9444 295576 9450
rect 295524 9386 295576 9392
rect 295996 6322 296024 335650
rect 296444 335640 296496 335646
rect 296444 335582 296496 335588
rect 296456 333946 296484 335582
rect 296548 334558 296576 336602
rect 296628 336592 296680 336598
rect 296628 336534 296680 336540
rect 296536 334552 296588 334558
rect 296536 334494 296588 334500
rect 296444 333940 296496 333946
rect 296444 333882 296496 333888
rect 295984 6316 296036 6322
rect 295984 6258 296036 6264
rect 294236 5704 294288 5710
rect 294236 5646 294288 5652
rect 288992 4344 289044 4350
rect 288992 4286 289044 4292
rect 287796 3392 287848 3398
rect 287796 3334 287848 3340
rect 288348 3392 288400 3398
rect 288348 3334 288400 3340
rect 287808 480 287836 3334
rect 289004 480 289032 4286
rect 292580 4276 292632 4282
rect 292580 4218 292632 4224
rect 291384 3732 291436 3738
rect 291384 3674 291436 3680
rect 290186 3632 290242 3641
rect 290186 3567 290242 3576
rect 290200 480 290228 3567
rect 291396 480 291424 3674
rect 292592 480 292620 4218
rect 293684 3800 293736 3806
rect 293684 3742 293736 3748
rect 294878 3768 294934 3777
rect 293696 480 293724 3742
rect 294878 3703 294934 3712
rect 294892 480 294920 3703
rect 296640 3398 296668 336534
rect 296732 336530 296760 338014
rect 296916 336666 296944 338014
rect 296904 336660 296956 336666
rect 296904 336602 296956 336608
rect 296720 336524 296772 336530
rect 296720 336466 296772 336472
rect 297284 335354 297312 338014
rect 296824 335326 297312 335354
rect 296824 9518 296852 335326
rect 297652 316034 297680 338014
rect 298112 335646 298140 338014
rect 298100 335640 298152 335646
rect 298100 335582 298152 335588
rect 298388 335354 298416 338014
rect 296916 316006 297680 316034
rect 298204 335326 298416 335354
rect 296812 9512 296864 9518
rect 296812 9454 296864 9460
rect 296916 5234 296944 316006
rect 298204 9586 298232 335326
rect 298756 316034 298784 338014
rect 299124 333198 299152 338014
rect 299388 336524 299440 336530
rect 299388 336466 299440 336472
rect 299112 333192 299164 333198
rect 299112 333134 299164 333140
rect 298296 316006 298784 316034
rect 298192 9580 298244 9586
rect 298192 9522 298244 9528
rect 298296 5302 298324 316006
rect 298284 5296 298336 5302
rect 298284 5238 298336 5244
rect 296904 5228 296956 5234
rect 296904 5170 296956 5176
rect 297272 3868 297324 3874
rect 297272 3810 297324 3816
rect 296076 3392 296128 3398
rect 296076 3334 296128 3340
rect 296628 3392 296680 3398
rect 296628 3334 296680 3340
rect 296088 480 296116 3334
rect 297284 480 297312 3810
rect 299400 3398 299428 336466
rect 299572 330064 299624 330070
rect 299572 330006 299624 330012
rect 299584 8906 299612 330006
rect 299676 9654 299704 338014
rect 299860 316034 299888 338014
rect 300228 335850 300256 338014
rect 300492 336728 300544 336734
rect 300492 336670 300544 336676
rect 300216 335844 300268 335850
rect 300216 335786 300268 335792
rect 300504 334490 300532 336670
rect 300492 334484 300544 334490
rect 300492 334426 300544 334432
rect 300596 330070 300624 338014
rect 300768 336660 300820 336666
rect 300768 336602 300820 336608
rect 300584 330064 300636 330070
rect 300584 330006 300636 330012
rect 299768 316006 299888 316034
rect 299664 9648 299716 9654
rect 299664 9590 299716 9596
rect 299572 8900 299624 8906
rect 299572 8842 299624 8848
rect 299664 6384 299716 6390
rect 299664 6326 299716 6332
rect 298468 3392 298520 3398
rect 298468 3334 298520 3340
rect 299388 3392 299440 3398
rect 299388 3334 299440 3340
rect 298480 480 298508 3334
rect 299676 480 299704 6326
rect 299768 5370 299796 316006
rect 299756 5364 299808 5370
rect 299756 5306 299808 5312
rect 300780 480 300808 336602
rect 300952 330540 301004 330546
rect 300952 330482 301004 330488
rect 300964 8838 300992 330482
rect 300952 8832 301004 8838
rect 300952 8774 301004 8780
rect 301056 5438 301084 338014
rect 301332 336734 301360 338014
rect 301320 336728 301372 336734
rect 301320 336670 301372 336676
rect 301700 330546 301728 338014
rect 302298 337770 302326 338028
rect 302436 338014 302680 338042
rect 302804 338014 303048 338042
rect 303172 338014 303416 338042
rect 303632 338014 303784 338042
rect 303908 338014 304152 338042
rect 304276 338014 304520 338042
rect 304644 338014 304888 338042
rect 305196 338014 305256 338042
rect 305380 338014 305624 338042
rect 305748 338014 305992 338042
rect 306116 338014 306360 338042
rect 306484 338014 306728 338042
rect 306852 338014 307096 338042
rect 307220 338014 307372 338042
rect 307496 338014 307740 338042
rect 307864 338014 308108 338042
rect 308232 338014 308476 338042
rect 308600 338014 308844 338042
rect 302298 337742 302372 337770
rect 301688 330540 301740 330546
rect 301688 330482 301740 330488
rect 302344 5506 302372 337742
rect 302436 332586 302464 338014
rect 302804 335354 302832 338014
rect 302528 335326 302832 335354
rect 302424 332580 302476 332586
rect 302424 332522 302476 332528
rect 302528 330562 302556 335326
rect 302436 330534 302556 330562
rect 302436 8770 302464 330534
rect 303172 316034 303200 338014
rect 303632 334422 303660 338014
rect 303908 335354 303936 338014
rect 303724 335326 303936 335354
rect 303620 334416 303672 334422
rect 303620 334358 303672 334364
rect 302528 316006 303200 316034
rect 302424 8764 302476 8770
rect 302424 8706 302476 8712
rect 302332 5500 302384 5506
rect 302332 5442 302384 5448
rect 301044 5432 301096 5438
rect 301044 5374 301096 5380
rect 302528 4758 302556 316006
rect 303724 8702 303752 335326
rect 304276 316034 304304 338014
rect 304644 333130 304672 338014
rect 304908 336728 304960 336734
rect 304908 336670 304960 336676
rect 304632 333124 304684 333130
rect 304632 333066 304684 333072
rect 303816 316006 304304 316034
rect 303712 8696 303764 8702
rect 303712 8638 303764 8644
rect 303160 6316 303212 6322
rect 303160 6258 303212 6264
rect 302516 4752 302568 4758
rect 302516 4694 302568 4700
rect 301964 3936 302016 3942
rect 301964 3878 302016 3884
rect 301976 480 302004 3878
rect 303172 480 303200 6258
rect 303816 4690 303844 316006
rect 303804 4684 303856 4690
rect 303804 4626 303856 4632
rect 304920 2990 304948 336670
rect 305196 330562 305224 338014
rect 305092 330540 305144 330546
rect 305196 330534 305316 330562
rect 305092 330482 305144 330488
rect 305000 326936 305052 326942
rect 305000 326878 305052 326884
rect 305012 4622 305040 326878
rect 305104 7138 305132 330482
rect 305184 330472 305236 330478
rect 305184 330414 305236 330420
rect 305196 8566 305224 330414
rect 305288 8634 305316 330534
rect 305380 326942 305408 338014
rect 305748 330546 305776 338014
rect 305736 330540 305788 330546
rect 305736 330482 305788 330488
rect 306116 330478 306144 338014
rect 306484 335354 306512 338014
rect 306852 335354 306880 338014
rect 306392 335326 306512 335354
rect 306576 335326 306880 335354
rect 306104 330472 306156 330478
rect 306104 330414 306156 330420
rect 305368 326936 305420 326942
rect 305368 326878 305420 326884
rect 305276 8628 305328 8634
rect 305276 8570 305328 8576
rect 305184 8560 305236 8566
rect 305184 8502 305236 8508
rect 305092 7132 305144 7138
rect 305092 7074 305144 7080
rect 305000 4616 305052 4622
rect 305000 4558 305052 4564
rect 306392 4554 306420 335326
rect 306472 326528 306524 326534
rect 306472 326470 306524 326476
rect 306484 4826 306512 326470
rect 306576 7070 306604 335326
rect 307220 316034 307248 338014
rect 307496 326534 307524 338014
rect 307760 330540 307812 330546
rect 307760 330482 307812 330488
rect 307484 326528 307536 326534
rect 307484 326470 307536 326476
rect 306668 316006 307248 316034
rect 306668 8498 306696 316006
rect 306656 8492 306708 8498
rect 306656 8434 306708 8440
rect 306564 7064 306616 7070
rect 306564 7006 306616 7012
rect 307772 4894 307800 330482
rect 307864 7614 307892 338014
rect 308232 316034 308260 338014
rect 308600 330546 308628 338014
rect 309198 337770 309226 338028
rect 309428 338014 309580 338042
rect 309704 338014 309948 338042
rect 310072 338014 310316 338042
rect 309198 337742 309272 337770
rect 308588 330540 308640 330546
rect 308588 330482 308640 330488
rect 309140 330472 309192 330478
rect 309140 330414 309192 330420
rect 307956 316006 308260 316034
rect 307956 8974 307984 316006
rect 307944 8968 307996 8974
rect 307944 8910 307996 8916
rect 307852 7608 307904 7614
rect 307852 7550 307904 7556
rect 309152 4962 309180 330414
rect 309244 7682 309272 337742
rect 309324 330540 309376 330546
rect 309324 330482 309376 330488
rect 309336 7750 309364 330482
rect 309428 8430 309456 338014
rect 309704 330478 309732 338014
rect 310072 330546 310100 338014
rect 310670 337770 310698 338028
rect 310808 338014 311052 338042
rect 311176 338014 311420 338042
rect 311544 338014 311788 338042
rect 311912 338014 312156 338042
rect 312280 338014 312524 338042
rect 312648 338014 312892 338042
rect 313016 338014 313260 338042
rect 313384 338014 313628 338042
rect 313752 338014 313996 338042
rect 314120 338014 314364 338042
rect 314732 338014 314884 338042
rect 310670 337742 310744 337770
rect 310520 336796 310572 336802
rect 310520 336738 310572 336744
rect 310060 330540 310112 330546
rect 310060 330482 310112 330488
rect 309692 330472 309744 330478
rect 309692 330414 309744 330420
rect 309416 8424 309468 8430
rect 309416 8366 309468 8372
rect 309324 7744 309376 7750
rect 309324 7686 309376 7692
rect 309232 7676 309284 7682
rect 309232 7618 309284 7624
rect 310532 5030 310560 336738
rect 310612 330540 310664 330546
rect 310612 330482 310664 330488
rect 310624 7818 310652 330482
rect 310716 9042 310744 337742
rect 310808 336802 310836 338014
rect 310796 336796 310848 336802
rect 310796 336738 310848 336744
rect 311176 330546 311204 338014
rect 311164 330540 311216 330546
rect 311164 330482 311216 330488
rect 311544 316034 311572 338014
rect 311912 335918 311940 338014
rect 311900 335912 311952 335918
rect 311900 335854 311952 335860
rect 311992 330540 312044 330546
rect 311992 330482 312044 330488
rect 310808 316006 311572 316034
rect 310808 9110 310836 316006
rect 312004 14482 312032 330482
rect 312280 316034 312308 338014
rect 312648 330546 312676 338014
rect 313016 335782 313044 338014
rect 313004 335776 313056 335782
rect 313004 335718 313056 335724
rect 312636 330540 312688 330546
rect 312636 330482 312688 330488
rect 313280 330540 313332 330546
rect 313280 330482 313332 330488
rect 312096 316006 312308 316034
rect 311992 14476 312044 14482
rect 311992 14418 312044 14424
rect 310796 9104 310848 9110
rect 310796 9046 310848 9052
rect 310704 9036 310756 9042
rect 310704 8978 310756 8984
rect 312096 7886 312124 316006
rect 312084 7880 312136 7886
rect 312084 7822 312136 7828
rect 310612 7812 310664 7818
rect 310612 7754 310664 7760
rect 313292 6186 313320 330482
rect 313384 7954 313412 338014
rect 313752 316034 313780 338014
rect 314120 330546 314148 338014
rect 314108 330540 314160 330546
rect 314108 330482 314160 330488
rect 314752 327208 314804 327214
rect 314752 327150 314804 327156
rect 313476 316006 313780 316034
rect 313476 10334 313504 316006
rect 313464 10328 313516 10334
rect 313464 10270 313516 10276
rect 314764 8090 314792 327150
rect 314752 8084 314804 8090
rect 314752 8026 314804 8032
rect 314856 8022 314884 338014
rect 314948 338014 315100 338042
rect 315224 338014 315468 338042
rect 315592 338014 315836 338042
rect 316052 338014 316204 338042
rect 316328 338014 316572 338042
rect 316696 338014 316940 338042
rect 317064 338014 317308 338042
rect 317524 338014 317676 338042
rect 317800 338014 318044 338042
rect 318168 338014 318412 338042
rect 318536 338014 318780 338042
rect 318996 338014 319148 338042
rect 319272 338014 319424 338042
rect 319548 338014 319792 338042
rect 319916 338014 320160 338042
rect 320284 338014 320528 338042
rect 320652 338014 320896 338042
rect 321020 338014 321264 338042
rect 321572 338014 321632 338042
rect 321756 338014 322000 338042
rect 322124 338014 322368 338042
rect 322492 338014 322736 338042
rect 323044 338014 323104 338042
rect 323228 338014 323472 338042
rect 323596 338014 323840 338042
rect 323964 338014 324208 338042
rect 324424 338014 324576 338042
rect 324700 338014 324944 338042
rect 325068 338014 325312 338042
rect 325436 338014 325680 338042
rect 325988 338014 326048 338042
rect 326172 338014 326416 338042
rect 326540 338014 326784 338042
rect 327092 338014 327152 338042
rect 327276 338014 327520 338042
rect 327644 338014 327888 338042
rect 328012 338014 328256 338042
rect 328472 338014 328624 338042
rect 328748 338014 328992 338042
rect 329116 338014 329360 338042
rect 329484 338014 329728 338042
rect 329852 338014 330096 338042
rect 330220 338014 330464 338042
rect 330588 338014 330832 338042
rect 330956 338014 331108 338042
rect 331416 338014 331476 338042
rect 331600 338014 331844 338042
rect 331968 338014 332212 338042
rect 332336 338014 332580 338042
rect 332796 338014 332948 338042
rect 333072 338014 333316 338042
rect 333440 338014 333684 338042
rect 333992 338014 334052 338042
rect 334360 338014 334420 338042
rect 334544 338014 334788 338042
rect 334912 338014 335156 338042
rect 335464 338014 335524 338042
rect 335648 338014 335892 338042
rect 336016 338014 336260 338042
rect 336384 338014 336628 338042
rect 336752 338014 336996 338042
rect 337120 338014 337364 338042
rect 337488 338014 337732 338042
rect 337856 338014 338100 338042
rect 338224 338014 338468 338042
rect 338592 338014 338836 338042
rect 338960 338014 339204 338042
rect 314948 335714 314976 338014
rect 315224 335986 315252 338014
rect 315212 335980 315264 335986
rect 315212 335922 315264 335928
rect 314936 335708 314988 335714
rect 314936 335650 314988 335656
rect 315592 327214 315620 338014
rect 316052 336054 316080 338014
rect 316328 336682 316356 338014
rect 316144 336654 316356 336682
rect 316040 336048 316092 336054
rect 316040 335990 316092 335996
rect 315580 327208 315632 327214
rect 315580 327150 315632 327156
rect 316144 10402 316172 336654
rect 316696 336546 316724 338014
rect 316236 336518 316724 336546
rect 316132 10396 316184 10402
rect 316132 10338 316184 10344
rect 316236 8158 316264 336518
rect 317064 336190 317092 338014
rect 317052 336184 317104 336190
rect 317052 336126 317104 336132
rect 316684 336048 316736 336054
rect 316684 335990 316736 335996
rect 316224 8152 316276 8158
rect 316224 8094 316276 8100
rect 314844 8016 314896 8022
rect 314844 7958 314896 7964
rect 313372 7948 313424 7954
rect 313372 7890 313424 7896
rect 316696 6390 316724 335990
rect 317524 10470 317552 338014
rect 317604 330540 317656 330546
rect 317604 330482 317656 330488
rect 317616 10538 317644 330482
rect 317800 316034 317828 338014
rect 318168 336122 318196 338014
rect 318156 336116 318208 336122
rect 318156 336058 318208 336064
rect 318536 330546 318564 338014
rect 318524 330540 318576 330546
rect 318524 330482 318576 330488
rect 318892 330540 318944 330546
rect 318892 330482 318944 330488
rect 317708 316006 317828 316034
rect 317604 10532 317656 10538
rect 317604 10474 317656 10480
rect 317512 10464 317564 10470
rect 317512 10406 317564 10412
rect 316684 6384 316736 6390
rect 316684 6326 316736 6332
rect 317708 6254 317736 316006
rect 317696 6248 317748 6254
rect 317696 6190 317748 6196
rect 313280 6180 313332 6186
rect 313280 6122 313332 6128
rect 318904 5098 318932 330482
rect 318892 5092 318944 5098
rect 318892 5034 318944 5040
rect 310520 5024 310572 5030
rect 310520 4966 310572 4972
rect 309140 4956 309192 4962
rect 309140 4898 309192 4904
rect 307760 4888 307812 4894
rect 307760 4830 307812 4836
rect 306472 4820 306524 4826
rect 306472 4762 306524 4768
rect 306380 4548 306432 4554
rect 306380 4490 306432 4496
rect 306748 4140 306800 4146
rect 306748 4082 306800 4088
rect 305552 4004 305604 4010
rect 305552 3946 305604 3952
rect 304356 2984 304408 2990
rect 304356 2926 304408 2932
rect 304908 2984 304960 2990
rect 304908 2926 304960 2932
rect 304368 480 304396 2926
rect 305564 480 305592 3946
rect 306760 480 306788 4082
rect 309048 4072 309100 4078
rect 309048 4014 309100 4020
rect 307944 3392 307996 3398
rect 307944 3334 307996 3340
rect 307956 480 307984 3334
rect 309060 480 309088 4014
rect 318996 3466 319024 338014
rect 319272 336258 319300 338014
rect 319260 336252 319312 336258
rect 319260 336194 319312 336200
rect 319548 330546 319576 338014
rect 319916 336394 319944 338014
rect 319904 336388 319956 336394
rect 319904 336330 319956 336336
rect 320284 335354 320312 338014
rect 320192 335326 320312 335354
rect 319536 330540 319588 330546
rect 319536 330482 319588 330488
rect 318984 3460 319036 3466
rect 318984 3402 319036 3408
rect 319720 3460 319772 3466
rect 319720 3402 319772 3408
rect 310244 3324 310296 3330
rect 310244 3266 310296 3272
rect 310256 480 310284 3266
rect 312636 3256 312688 3262
rect 312636 3198 312688 3204
rect 311440 3188 311492 3194
rect 311440 3130 311492 3136
rect 311452 480 311480 3130
rect 312648 480 312676 3198
rect 313832 3120 313884 3126
rect 313832 3062 313884 3068
rect 313844 480 313872 3062
rect 317328 3052 317380 3058
rect 317328 2994 317380 3000
rect 315028 2984 315080 2990
rect 315028 2926 315080 2932
rect 315040 480 315068 2926
rect 316224 2916 316276 2922
rect 316224 2858 316276 2864
rect 316236 480 316264 2858
rect 317340 480 317368 2994
rect 318524 2848 318576 2854
rect 318524 2790 318576 2796
rect 318536 480 318564 2790
rect 319732 480 319760 3402
rect 320192 3369 320220 335326
rect 320272 330540 320324 330546
rect 320272 330482 320324 330488
rect 320284 3534 320312 330482
rect 320652 316034 320680 338014
rect 321020 330546 321048 338014
rect 321572 336326 321600 338014
rect 321560 336320 321612 336326
rect 321560 336262 321612 336268
rect 321008 330540 321060 330546
rect 321008 330482 321060 330488
rect 321652 330540 321704 330546
rect 321652 330482 321704 330488
rect 320376 316006 320680 316034
rect 320376 5166 320404 316006
rect 320364 5160 320416 5166
rect 320364 5102 320416 5108
rect 320916 3868 320968 3874
rect 320916 3810 320968 3816
rect 320272 3528 320324 3534
rect 320272 3470 320324 3476
rect 320178 3360 320234 3369
rect 320178 3295 320234 3304
rect 320928 480 320956 3810
rect 321664 3505 321692 330482
rect 321756 4486 321784 338014
rect 322124 330546 322152 338014
rect 322112 330540 322164 330546
rect 322112 330482 322164 330488
rect 322492 316034 322520 338014
rect 321848 316006 322520 316034
rect 321744 4480 321796 4486
rect 321744 4422 321796 4428
rect 321848 3670 321876 316006
rect 323044 4418 323072 338014
rect 323124 330540 323176 330546
rect 323124 330482 323176 330488
rect 323032 4412 323084 4418
rect 323032 4354 323084 4360
rect 323136 4350 323164 330482
rect 323124 4344 323176 4350
rect 323124 4286 323176 4292
rect 321836 3664 321888 3670
rect 321836 3606 321888 3612
rect 323228 3602 323256 338014
rect 323596 336462 323624 338014
rect 323584 336456 323636 336462
rect 323584 336398 323636 336404
rect 323964 330546 323992 338014
rect 324424 330818 324452 338014
rect 324700 335354 324728 338014
rect 324516 335326 324728 335354
rect 324412 330812 324464 330818
rect 324412 330754 324464 330760
rect 324516 330698 324544 335326
rect 324332 330670 324544 330698
rect 323952 330540 324004 330546
rect 323952 330482 324004 330488
rect 324332 3738 324360 330670
rect 324412 330608 324464 330614
rect 324412 330550 324464 330556
rect 324424 3913 324452 330550
rect 324504 330540 324556 330546
rect 324504 330482 324556 330488
rect 324410 3904 324466 3913
rect 324410 3839 324466 3848
rect 324320 3732 324372 3738
rect 324320 3674 324372 3680
rect 324412 3732 324464 3738
rect 324412 3674 324464 3680
rect 323216 3596 323268 3602
rect 323216 3538 323268 3544
rect 323308 3596 323360 3602
rect 323308 3538 323360 3544
rect 322112 3528 322164 3534
rect 321650 3496 321706 3505
rect 322112 3470 322164 3476
rect 321650 3431 321706 3440
rect 322124 480 322152 3470
rect 323320 480 323348 3538
rect 324424 480 324452 3674
rect 324516 3670 324544 330482
rect 325068 316034 325096 338014
rect 325436 330546 325464 338014
rect 325424 330540 325476 330546
rect 325424 330482 325476 330488
rect 325792 330540 325844 330546
rect 325792 330482 325844 330488
rect 324608 316006 325096 316034
rect 324608 4282 324636 316006
rect 324596 4276 324648 4282
rect 324596 4218 324648 4224
rect 325804 3942 325832 330482
rect 325988 4049 326016 338014
rect 326172 336598 326200 338014
rect 326160 336592 326212 336598
rect 326160 336534 326212 336540
rect 326540 330546 326568 338014
rect 327092 336530 327120 338014
rect 327080 336524 327132 336530
rect 327080 336466 327132 336472
rect 327276 336054 327304 338014
rect 327644 336818 327672 338014
rect 327552 336790 327672 336818
rect 327552 336666 327580 336790
rect 328012 336682 328040 338014
rect 327540 336660 327592 336666
rect 327540 336602 327592 336608
rect 327644 336654 328040 336682
rect 327264 336048 327316 336054
rect 327264 335990 327316 335996
rect 326528 330540 326580 330546
rect 326528 330482 326580 330488
rect 327644 316034 327672 336654
rect 328472 336598 328500 338014
rect 328748 336734 328776 338014
rect 328736 336728 328788 336734
rect 328736 336670 328788 336676
rect 327724 336592 327776 336598
rect 327724 336534 327776 336540
rect 328460 336592 328512 336598
rect 328460 336534 328512 336540
rect 327276 316006 327672 316034
rect 325974 4040 326030 4049
rect 325974 3975 326030 3984
rect 325792 3936 325844 3942
rect 325792 3878 325844 3884
rect 326804 3936 326856 3942
rect 326804 3878 326856 3884
rect 324504 3664 324556 3670
rect 324504 3606 324556 3612
rect 325608 3664 325660 3670
rect 325608 3606 325660 3612
rect 325620 480 325648 3606
rect 326816 480 326844 3878
rect 327276 3806 327304 316006
rect 327736 6322 327764 336534
rect 328368 336116 328420 336122
rect 328368 336058 328420 336064
rect 328380 6914 328408 336058
rect 329116 335354 329144 338014
rect 329196 336728 329248 336734
rect 329196 336670 329248 336676
rect 329024 335326 329144 335354
rect 328552 330540 328604 330546
rect 328552 330482 328604 330488
rect 328012 6886 328408 6914
rect 327724 6316 327776 6322
rect 327724 6258 327776 6264
rect 327264 3800 327316 3806
rect 327264 3742 327316 3748
rect 328012 480 328040 6886
rect 328564 4146 328592 330482
rect 329024 316034 329052 335326
rect 329208 316034 329236 336670
rect 329484 330546 329512 338014
rect 329472 330540 329524 330546
rect 329472 330482 329524 330488
rect 328748 316006 329052 316034
rect 329116 316006 329236 316034
rect 328552 4140 328604 4146
rect 328552 4082 328604 4088
rect 328748 4010 328776 316006
rect 328736 4004 328788 4010
rect 328736 3946 328788 3952
rect 329116 3874 329144 316006
rect 329196 4004 329248 4010
rect 329196 3946 329248 3952
rect 329104 3868 329156 3874
rect 329104 3810 329156 3816
rect 329208 480 329236 3946
rect 329852 3398 329880 338014
rect 330024 330540 330076 330546
rect 330024 330482 330076 330488
rect 329932 330472 329984 330478
rect 329932 330414 329984 330420
rect 329840 3392 329892 3398
rect 329840 3334 329892 3340
rect 329944 3194 329972 330414
rect 330036 3330 330064 330482
rect 330220 316034 330248 338014
rect 330588 330546 330616 338014
rect 330576 330540 330628 330546
rect 330576 330482 330628 330488
rect 330956 330478 330984 338014
rect 331312 330540 331364 330546
rect 331312 330482 331364 330488
rect 330944 330472 330996 330478
rect 330944 330414 330996 330420
rect 330128 316006 330248 316034
rect 330128 4078 330156 316006
rect 330116 4072 330168 4078
rect 330116 4014 330168 4020
rect 330392 3460 330444 3466
rect 330392 3402 330444 3408
rect 330024 3324 330076 3330
rect 330024 3266 330076 3272
rect 329932 3188 329984 3194
rect 329932 3130 329984 3136
rect 330404 480 330432 3402
rect 331324 2922 331352 330482
rect 331416 3262 331444 338014
rect 331600 335354 331628 338014
rect 331508 335326 331628 335354
rect 331404 3256 331456 3262
rect 331404 3198 331456 3204
rect 331508 3126 331536 335326
rect 331968 316034 331996 338014
rect 332336 330546 332364 338014
rect 332508 335368 332560 335374
rect 332508 335310 332560 335316
rect 332324 330540 332376 330546
rect 332324 330482 332376 330488
rect 331600 316006 331996 316034
rect 331600 16574 331628 316006
rect 331600 16546 331720 16574
rect 331588 3528 331640 3534
rect 331588 3470 331640 3476
rect 331496 3120 331548 3126
rect 331496 3062 331548 3068
rect 331312 2916 331364 2922
rect 331312 2858 331364 2864
rect 331600 480 331628 3470
rect 331692 2990 331720 16546
rect 332520 3534 332548 335310
rect 332692 330540 332744 330546
rect 332692 330482 332744 330488
rect 332600 330200 332652 330206
rect 332600 330142 332652 330148
rect 332612 4282 332640 330142
rect 332600 4276 332652 4282
rect 332600 4218 332652 4224
rect 332704 4162 332732 330482
rect 332796 16574 332824 338014
rect 333072 330206 333100 338014
rect 333244 336048 333296 336054
rect 333244 335990 333296 335996
rect 333060 330200 333112 330206
rect 333060 330142 333112 330148
rect 332796 16546 333008 16574
rect 332784 4276 332836 4282
rect 332784 4218 332836 4224
rect 332612 4134 332732 4162
rect 332612 3602 332640 4134
rect 332692 4072 332744 4078
rect 332692 4014 332744 4020
rect 332600 3596 332652 3602
rect 332600 3538 332652 3544
rect 332508 3528 332560 3534
rect 332508 3470 332560 3476
rect 331680 2984 331732 2990
rect 331680 2926 331732 2932
rect 332704 480 332732 4014
rect 332796 2854 332824 4218
rect 332980 3058 333008 16546
rect 333256 3466 333284 335990
rect 333440 330546 333468 338014
rect 333992 336734 334020 338014
rect 333980 336728 334032 336734
rect 333980 336670 334032 336676
rect 333428 330540 333480 330546
rect 333428 330482 333480 330488
rect 334072 330540 334124 330546
rect 334072 330482 334124 330488
rect 333888 3868 333940 3874
rect 333888 3810 333940 3816
rect 333244 3460 333296 3466
rect 333244 3402 333296 3408
rect 332968 3052 333020 3058
rect 332968 2994 333020 3000
rect 332784 2848 332836 2854
rect 332784 2790 332836 2796
rect 333900 480 333928 3810
rect 334084 3806 334112 330482
rect 334164 326732 334216 326738
rect 334164 326674 334216 326680
rect 334072 3800 334124 3806
rect 334072 3742 334124 3748
rect 334176 3738 334204 326674
rect 334164 3732 334216 3738
rect 334164 3674 334216 3680
rect 334360 3398 334388 338014
rect 334544 330546 334572 338014
rect 334532 330540 334584 330546
rect 334532 330482 334584 330488
rect 334912 326738 334940 338014
rect 334900 326732 334952 326738
rect 334900 326674 334952 326680
rect 335464 3670 335492 338014
rect 335544 330540 335596 330546
rect 335544 330482 335596 330488
rect 335556 4010 335584 330482
rect 335544 4004 335596 4010
rect 335544 3946 335596 3952
rect 335648 3942 335676 338014
rect 336016 336122 336044 338014
rect 336004 336116 336056 336122
rect 336004 336058 336056 336064
rect 336004 335980 336056 335986
rect 336004 335922 336056 335928
rect 336016 4078 336044 335922
rect 336384 330546 336412 338014
rect 336752 336054 336780 338014
rect 336740 336048 336792 336054
rect 336740 335990 336792 335996
rect 337120 335374 337148 338014
rect 337488 335986 337516 338014
rect 337476 335980 337528 335986
rect 337476 335922 337528 335928
rect 337108 335368 337160 335374
rect 337108 335310 337160 335316
rect 336372 330540 336424 330546
rect 336372 330482 336424 330488
rect 337856 316034 337884 338014
rect 338120 330540 338172 330546
rect 338120 330482 338172 330488
rect 336936 316006 337884 316034
rect 336004 4072 336056 4078
rect 336004 4014 336056 4020
rect 335636 3936 335688 3942
rect 335636 3878 335688 3884
rect 336936 3874 336964 316006
rect 336924 3868 336976 3874
rect 336924 3810 336976 3816
rect 335452 3664 335504 3670
rect 335452 3606 335504 3612
rect 338132 3534 338160 330482
rect 337476 3528 337528 3534
rect 337476 3470 337528 3476
rect 338120 3528 338172 3534
rect 338120 3470 338172 3476
rect 335084 3460 335136 3466
rect 335084 3402 335136 3408
rect 334348 3392 334400 3398
rect 334348 3334 334400 3340
rect 335096 480 335124 3402
rect 336280 2984 336332 2990
rect 336280 2926 336332 2932
rect 336292 480 336320 2926
rect 337488 480 337516 3470
rect 338224 3466 338252 338014
rect 338592 316034 338620 338014
rect 338960 330546 338988 338014
rect 339558 337770 339586 338028
rect 339788 338014 339940 338042
rect 340308 338014 340552 338042
rect 340676 338014 340828 338042
rect 341044 338014 341288 338042
rect 341412 338014 341656 338042
rect 341780 338014 342024 338042
rect 339558 337742 339632 337770
rect 339500 336728 339552 336734
rect 339500 336670 339552 336676
rect 338948 330540 339000 330546
rect 338948 330482 339000 330488
rect 338316 316006 338620 316034
rect 338212 3460 338264 3466
rect 338212 3402 338264 3408
rect 338316 2990 338344 316006
rect 338672 3120 338724 3126
rect 338672 3062 338724 3068
rect 338304 2984 338356 2990
rect 338304 2926 338356 2932
rect 338684 480 338712 3062
rect 339512 2938 339540 336670
rect 339604 3126 339632 337742
rect 339788 336734 339816 338014
rect 339776 336728 339828 336734
rect 339776 336670 339828 336676
rect 340524 335354 340552 338014
rect 340800 336682 340828 338014
rect 340800 336654 341196 336682
rect 340524 335326 340828 335354
rect 340800 3482 340828 335326
rect 341168 16574 341196 336654
rect 341260 335578 341288 338014
rect 341628 336734 341656 338014
rect 341616 336728 341668 336734
rect 341616 336670 341668 336676
rect 341248 335572 341300 335578
rect 341248 335514 341300 335520
rect 341996 335442 342024 338014
rect 342134 337770 342162 338028
rect 342516 338014 342760 338042
rect 342884 338014 343036 338042
rect 343160 338014 343404 338042
rect 342134 337742 342208 337770
rect 342076 336728 342128 336734
rect 342076 336670 342128 336676
rect 341984 335436 342036 335442
rect 341984 335378 342036 335384
rect 341168 16546 342024 16574
rect 341996 3482 342024 16546
rect 342088 3602 342116 336670
rect 342180 4010 342208 337742
rect 342732 335714 342760 338014
rect 342720 335708 342772 335714
rect 342720 335650 342772 335656
rect 342352 335572 342404 335578
rect 342352 335514 342404 335520
rect 342364 16574 342392 335514
rect 343008 325694 343036 338014
rect 343376 336682 343404 338014
rect 343514 337770 343542 338028
rect 343896 338014 344140 338042
rect 344264 338014 344508 338042
rect 344632 338014 344876 338042
rect 343514 337742 343588 337770
rect 343560 336734 343588 337742
rect 343548 336728 343600 336734
rect 343376 336654 343496 336682
rect 343548 336670 343600 336676
rect 343364 335708 343416 335714
rect 343364 335650 343416 335656
rect 343376 330426 343404 335650
rect 343468 330562 343496 336654
rect 344112 336190 344140 338014
rect 344284 336728 344336 336734
rect 344284 336670 344336 336676
rect 344100 336184 344152 336190
rect 344100 336126 344152 336132
rect 343468 330534 343588 330562
rect 343376 330398 343496 330426
rect 343008 325666 343404 325694
rect 342364 16546 343312 16574
rect 342168 4004 342220 4010
rect 342168 3946 342220 3952
rect 342076 3596 342128 3602
rect 342076 3538 342128 3544
rect 343284 3482 343312 16546
rect 343376 3806 343404 325666
rect 343468 4078 343496 330398
rect 343560 4146 343588 330534
rect 343548 4140 343600 4146
rect 343548 4082 343600 4088
rect 343456 4072 343508 4078
rect 343456 4014 343508 4020
rect 344296 3942 344324 336670
rect 344480 335510 344508 338014
rect 344848 336054 344876 338014
rect 344940 338014 345000 338042
rect 345368 338014 345612 338042
rect 345736 338014 345980 338042
rect 346104 338014 346348 338042
rect 346472 338014 346716 338042
rect 346840 338014 347084 338042
rect 347208 338014 347452 338042
rect 344836 336048 344888 336054
rect 344836 335990 344888 335996
rect 344468 335504 344520 335510
rect 344468 335446 344520 335452
rect 344940 335374 344968 338014
rect 345584 335850 345612 338014
rect 345664 336184 345716 336190
rect 345664 336126 345716 336132
rect 345572 335844 345624 335850
rect 345572 335786 345624 335792
rect 345112 335436 345164 335442
rect 345112 335378 345164 335384
rect 344928 335368 344980 335374
rect 344928 335310 344980 335316
rect 345124 16574 345152 335378
rect 345124 16546 345612 16574
rect 344284 3936 344336 3942
rect 344284 3878 344336 3884
rect 343364 3800 343416 3806
rect 343364 3742 343416 3748
rect 344560 3596 344612 3602
rect 344560 3538 344612 3544
rect 340800 3454 341012 3482
rect 341996 3454 342208 3482
rect 343284 3454 343404 3482
rect 339592 3120 339644 3126
rect 339592 3062 339644 3068
rect 339512 2910 339908 2938
rect 339880 480 339908 2910
rect 340984 480 341012 3454
rect 342180 480 342208 3454
rect 343376 480 343404 3454
rect 344572 480 344600 3538
rect 345584 3346 345612 16546
rect 345676 3534 345704 336126
rect 345756 335368 345808 335374
rect 345952 335354 345980 338014
rect 346320 336326 346348 338014
rect 346688 336394 346716 338014
rect 347056 336734 347084 338014
rect 347044 336728 347096 336734
rect 347044 336670 347096 336676
rect 347424 336530 347452 338014
rect 347516 338014 347576 338042
rect 347944 338014 348188 338042
rect 348312 338014 348464 338042
rect 348680 338014 348924 338042
rect 347412 336524 347464 336530
rect 347412 336466 347464 336472
rect 346676 336388 346728 336394
rect 346676 336330 346728 336336
rect 346308 336320 346360 336326
rect 346308 336262 346360 336268
rect 347136 336320 347188 336326
rect 347136 336262 347188 336268
rect 346952 335504 347004 335510
rect 346952 335446 347004 335452
rect 345952 335326 346348 335354
rect 345756 335310 345808 335316
rect 345768 3874 345796 335310
rect 345756 3868 345808 3874
rect 345756 3810 345808 3816
rect 346320 3738 346348 335326
rect 346964 325694 346992 335446
rect 346964 325666 347084 325694
rect 346952 4004 347004 4010
rect 346952 3946 347004 3952
rect 346308 3732 346360 3738
rect 346308 3674 346360 3680
rect 345664 3528 345716 3534
rect 345664 3470 345716 3476
rect 345584 3318 345796 3346
rect 345768 480 345796 3318
rect 346964 480 346992 3946
rect 347056 3126 347084 325666
rect 347148 3670 347176 336262
rect 347516 335578 347544 338014
rect 348160 336734 348188 338014
rect 347688 336728 347740 336734
rect 347688 336670 347740 336676
rect 348148 336728 348200 336734
rect 348148 336670 348200 336676
rect 347596 336388 347648 336394
rect 347596 336330 347648 336336
rect 347504 335572 347556 335578
rect 347504 335514 347556 335520
rect 347136 3664 347188 3670
rect 347136 3606 347188 3612
rect 347608 3602 347636 336330
rect 347596 3596 347648 3602
rect 347596 3538 347648 3544
rect 347700 3466 347728 336670
rect 348436 336598 348464 338014
rect 348424 336592 348476 336598
rect 348424 336534 348476 336540
rect 348896 336326 348924 338014
rect 348988 338014 349048 338042
rect 349416 338014 349660 338042
rect 349784 338014 350028 338042
rect 348884 336320 348936 336326
rect 348884 336262 348936 336268
rect 348424 336048 348476 336054
rect 348424 335990 348476 335996
rect 348056 4072 348108 4078
rect 348056 4014 348108 4020
rect 347688 3460 347740 3466
rect 347688 3402 347740 3408
rect 347044 3120 347096 3126
rect 347044 3062 347096 3068
rect 348068 480 348096 4014
rect 348436 3058 348464 335990
rect 348516 335572 348568 335578
rect 348516 335514 348568 335520
rect 348424 3052 348476 3058
rect 348424 2994 348476 3000
rect 348528 2990 348556 335514
rect 348988 3330 349016 338014
rect 349068 336728 349120 336734
rect 349068 336670 349120 336676
rect 348976 3324 349028 3330
rect 348976 3266 349028 3272
rect 349080 3262 349108 336670
rect 349632 335714 349660 338014
rect 349804 335844 349856 335850
rect 349804 335786 349856 335792
rect 349620 335708 349672 335714
rect 349620 335650 349672 335656
rect 349252 3800 349304 3806
rect 349252 3742 349304 3748
rect 349068 3256 349120 3262
rect 349068 3198 349120 3204
rect 348516 2984 348568 2990
rect 348516 2926 348568 2932
rect 349264 480 349292 3742
rect 349816 3194 349844 335786
rect 350000 330546 350028 338014
rect 350092 338014 350152 338042
rect 350276 338014 350520 338042
rect 350888 338014 351132 338042
rect 351256 338014 351500 338042
rect 351624 338014 351776 338042
rect 351992 338014 352236 338042
rect 352360 338014 352604 338042
rect 352728 338014 352880 338042
rect 350092 335442 350120 338014
rect 350080 335436 350132 335442
rect 350080 335378 350132 335384
rect 349988 330540 350040 330546
rect 349988 330482 350040 330488
rect 350276 4486 350304 338014
rect 351104 336734 351132 338014
rect 351092 336728 351144 336734
rect 351092 336670 351144 336676
rect 351472 336190 351500 338014
rect 351460 336184 351512 336190
rect 351460 336126 351512 336132
rect 350356 335436 350408 335442
rect 350356 335378 350408 335384
rect 350264 4480 350316 4486
rect 350264 4422 350316 4428
rect 350368 4078 350396 335378
rect 350448 330540 350500 330546
rect 350448 330482 350500 330488
rect 350460 4298 350488 330482
rect 351748 4554 351776 338014
rect 351828 336728 351880 336734
rect 351828 336670 351880 336676
rect 351736 4548 351788 4554
rect 351736 4490 351788 4496
rect 350460 4270 350580 4298
rect 350448 4140 350500 4146
rect 350448 4082 350500 4088
rect 350356 4072 350408 4078
rect 350356 4014 350408 4020
rect 349804 3188 349856 3194
rect 349804 3130 349856 3136
rect 350460 480 350488 4082
rect 350552 3398 350580 4270
rect 351840 4146 351868 336670
rect 352208 336462 352236 338014
rect 352196 336456 352248 336462
rect 352196 336398 352248 336404
rect 352576 335782 352604 338014
rect 352852 336734 352880 338014
rect 353036 338014 353096 338042
rect 353464 338014 353708 338042
rect 353832 338014 354076 338042
rect 354200 338014 354444 338042
rect 352840 336728 352892 336734
rect 352840 336670 352892 336676
rect 352564 335776 352616 335782
rect 352564 335718 352616 335724
rect 353036 10334 353064 338014
rect 353116 336728 353168 336734
rect 353116 336670 353168 336676
rect 353024 10328 353076 10334
rect 353024 10270 353076 10276
rect 353128 4622 353156 336670
rect 353680 336122 353708 338014
rect 354048 336258 354076 338014
rect 354416 336394 354444 338014
rect 354554 337770 354582 338028
rect 354936 338014 355088 338042
rect 355212 338014 355456 338042
rect 355580 338014 355732 338042
rect 354554 337742 354628 337770
rect 354404 336388 354456 336394
rect 354404 336330 354456 336336
rect 354036 336252 354088 336258
rect 354036 336194 354088 336200
rect 354496 336252 354548 336258
rect 354496 336194 354548 336200
rect 353668 336116 353720 336122
rect 353668 336058 353720 336064
rect 353208 335776 353260 335782
rect 353208 335718 353260 335724
rect 353116 4616 353168 4622
rect 353116 4558 353168 4564
rect 351828 4140 351880 4146
rect 351828 4082 351880 4088
rect 353220 4010 353248 335718
rect 353944 335708 353996 335714
rect 353944 335650 353996 335656
rect 353956 8974 353984 335650
rect 353944 8968 353996 8974
rect 353944 8910 353996 8916
rect 354508 4690 354536 336194
rect 354496 4684 354548 4690
rect 354496 4626 354548 4632
rect 353208 4004 353260 4010
rect 353208 3946 353260 3952
rect 354600 3942 354628 337742
rect 355060 336666 355088 338014
rect 355048 336660 355100 336666
rect 355048 336602 355100 336608
rect 355428 335374 355456 338014
rect 355704 336734 355732 338014
rect 355796 338014 355948 338042
rect 356316 338014 356560 338042
rect 356684 338014 356928 338042
rect 357052 338014 357296 338042
rect 355692 336728 355744 336734
rect 355692 336670 355744 336676
rect 355416 335368 355468 335374
rect 355416 335310 355468 335316
rect 355796 5506 355824 338014
rect 355968 336728 356020 336734
rect 355968 336670 356020 336676
rect 355876 336660 355928 336666
rect 355876 336602 355928 336608
rect 355784 5500 355836 5506
rect 355784 5442 355836 5448
rect 355888 4758 355916 336602
rect 355876 4752 355928 4758
rect 355876 4694 355928 4700
rect 351644 3936 351696 3942
rect 351644 3878 351696 3884
rect 354588 3936 354640 3942
rect 354588 3878 354640 3884
rect 350540 3392 350592 3398
rect 350540 3334 350592 3340
rect 351656 480 351684 3878
rect 355980 3806 356008 336670
rect 356532 336054 356560 338014
rect 356900 336598 356928 338014
rect 357164 336728 357216 336734
rect 357164 336670 357216 336676
rect 356888 336592 356940 336598
rect 356888 336534 356940 336540
rect 356520 336048 356572 336054
rect 356520 335990 356572 335996
rect 357176 9042 357204 336670
rect 357164 9036 357216 9042
rect 357164 8978 357216 8984
rect 357268 5438 357296 338014
rect 357360 338014 357420 338042
rect 357788 338014 358032 338042
rect 358156 338014 358400 338042
rect 357360 336734 357388 338014
rect 357348 336728 357400 336734
rect 357348 336670 357400 336676
rect 358004 336666 358032 338014
rect 358372 336734 358400 338014
rect 358510 337770 358538 338028
rect 358892 338014 359136 338042
rect 359260 338014 359504 338042
rect 359628 338014 359872 338042
rect 359996 338014 360148 338042
rect 360364 338014 360608 338042
rect 360732 338014 360976 338042
rect 361100 338014 361252 338042
rect 358510 337742 358584 337770
rect 358360 336728 358412 336734
rect 358360 336670 358412 336676
rect 357992 336660 358044 336666
rect 357992 336602 358044 336608
rect 357348 336592 357400 336598
rect 357348 336534 357400 336540
rect 357256 5432 357308 5438
rect 357256 5374 357308 5380
rect 357360 3874 357388 336534
rect 358084 336524 358136 336530
rect 358084 336466 358136 336472
rect 356336 3868 356388 3874
rect 356336 3810 356388 3816
rect 357348 3868 357400 3874
rect 357348 3810 357400 3816
rect 355968 3800 356020 3806
rect 355968 3742 356020 3748
rect 352840 3528 352892 3534
rect 352840 3470 352892 3476
rect 352852 480 352880 3470
rect 355232 3188 355284 3194
rect 355232 3130 355284 3136
rect 354036 3120 354088 3126
rect 354036 3062 354088 3068
rect 354048 480 354076 3062
rect 355244 480 355272 3130
rect 356348 480 356376 3810
rect 358096 3126 358124 336466
rect 358556 5370 358584 337742
rect 358636 336728 358688 336734
rect 358636 336670 358688 336676
rect 358544 5364 358596 5370
rect 358544 5306 358596 5312
rect 358648 5302 358676 336670
rect 358728 336660 358780 336666
rect 358728 336602 358780 336608
rect 358636 5296 358688 5302
rect 358636 5238 358688 5244
rect 358740 3806 358768 336602
rect 359108 335850 359136 338014
rect 359096 335844 359148 335850
rect 359096 335786 359148 335792
rect 359476 335354 359504 338014
rect 359844 336682 359872 338014
rect 359844 336654 359964 336682
rect 359476 335326 359872 335354
rect 359844 5234 359872 335326
rect 359832 5228 359884 5234
rect 359832 5170 359884 5176
rect 359936 5166 359964 336654
rect 360016 335844 360068 335850
rect 360016 335786 360068 335792
rect 359924 5160 359976 5166
rect 359924 5102 359976 5108
rect 358728 3800 358780 3806
rect 358728 3742 358780 3748
rect 360028 3670 360056 335786
rect 358728 3664 358780 3670
rect 358728 3606 358780 3612
rect 360016 3664 360068 3670
rect 360016 3606 360068 3612
rect 357532 3120 357584 3126
rect 357532 3062 357584 3068
rect 358084 3120 358136 3126
rect 358084 3062 358136 3068
rect 357544 480 357572 3062
rect 358740 480 358768 3606
rect 360120 3602 360148 338014
rect 360580 336734 360608 338014
rect 360568 336728 360620 336734
rect 360568 336670 360620 336676
rect 360948 326398 360976 338014
rect 361120 336728 361172 336734
rect 361120 336670 361172 336676
rect 360936 326392 360988 326398
rect 360936 326334 360988 326340
rect 361132 321554 361160 336670
rect 361224 335714 361252 338014
rect 361408 338014 361468 338042
rect 361836 338014 362080 338042
rect 362204 338014 362448 338042
rect 362572 338014 362816 338042
rect 361212 335708 361264 335714
rect 361212 335650 361264 335656
rect 361304 326392 361356 326398
rect 361304 326334 361356 326340
rect 361132 321526 361252 321554
rect 361224 5098 361252 321526
rect 361212 5092 361264 5098
rect 361212 5034 361264 5040
rect 361316 5030 361344 326334
rect 361304 5024 361356 5030
rect 361304 4966 361356 4972
rect 361408 4962 361436 338014
rect 362052 336666 362080 338014
rect 362040 336660 362092 336666
rect 362040 336602 362092 336608
rect 361488 335708 361540 335714
rect 361488 335650 361540 335656
rect 361396 4956 361448 4962
rect 361396 4898 361448 4904
rect 359924 3596 359976 3602
rect 359924 3538 359976 3544
rect 360108 3596 360160 3602
rect 360108 3538 360160 3544
rect 359936 480 359964 3538
rect 361500 3534 361528 335650
rect 362420 326398 362448 338014
rect 362592 336728 362644 336734
rect 362592 336670 362644 336676
rect 362408 326392 362460 326398
rect 362408 326334 362460 326340
rect 362604 7070 362632 336670
rect 362684 336660 362736 336666
rect 362684 336602 362736 336608
rect 362592 7064 362644 7070
rect 362592 7006 362644 7012
rect 362696 4894 362724 336602
rect 362684 4888 362736 4894
rect 362684 4830 362736 4836
rect 362788 4826 362816 338014
rect 362880 338014 362940 338042
rect 363308 338014 363552 338042
rect 363676 338014 363920 338042
rect 364044 338014 364196 338042
rect 364412 338014 364656 338042
rect 364780 338014 365024 338042
rect 365148 338014 365392 338042
rect 365516 338014 365668 338042
rect 365884 338014 366128 338042
rect 366252 338014 366496 338042
rect 366620 338014 366864 338042
rect 362880 336734 362908 338014
rect 363524 336734 363552 338014
rect 362868 336728 362920 336734
rect 362868 336670 362920 336676
rect 363512 336728 363564 336734
rect 363512 336670 363564 336676
rect 363604 336592 363656 336598
rect 363604 336534 363656 336540
rect 362868 326392 362920 326398
rect 362868 326334 362920 326340
rect 362776 4820 362828 4826
rect 362776 4762 362828 4768
rect 361120 3528 361172 3534
rect 361120 3470 361172 3476
rect 361488 3528 361540 3534
rect 361488 3470 361540 3476
rect 361132 480 361160 3470
rect 362880 3466 362908 326334
rect 363616 5574 363644 336534
rect 363892 335510 363920 338014
rect 363880 335504 363932 335510
rect 363880 335446 363932 335452
rect 364168 7138 364196 338014
rect 364248 336728 364300 336734
rect 364248 336670 364300 336676
rect 364156 7132 364208 7138
rect 364156 7074 364208 7080
rect 363604 5568 363656 5574
rect 363604 5510 363656 5516
rect 362316 3460 362368 3466
rect 362316 3402 362368 3408
rect 362868 3460 362920 3466
rect 362868 3402 362920 3408
rect 362328 480 362356 3402
rect 363512 3120 363564 3126
rect 363512 3062 363564 3068
rect 363524 480 363552 3062
rect 364260 2854 364288 336670
rect 364628 335442 364656 338014
rect 364996 335578 365024 338014
rect 364984 335572 365036 335578
rect 364984 335514 365036 335520
rect 364616 335436 364668 335442
rect 364616 335378 364668 335384
rect 365364 335354 365392 338014
rect 365364 335326 365576 335354
rect 365548 7206 365576 335326
rect 365536 7200 365588 7206
rect 365536 7142 365588 7148
rect 364616 3188 364668 3194
rect 364616 3130 364668 3136
rect 364248 2848 364300 2854
rect 364248 2790 364300 2796
rect 364628 480 364656 3130
rect 365640 2922 365668 338014
rect 366100 335646 366128 338014
rect 366468 336666 366496 338014
rect 366456 336660 366508 336666
rect 366456 336602 366508 336608
rect 366836 335714 366864 338014
rect 366928 338014 366988 338042
rect 367264 338014 367508 338042
rect 367632 338014 367876 338042
rect 368000 338014 368152 338042
rect 366928 335918 366956 338014
rect 367480 336734 367508 338014
rect 367468 336728 367520 336734
rect 367468 336670 367520 336676
rect 367008 336660 367060 336666
rect 367008 336602 367060 336608
rect 366916 335912 366968 335918
rect 366916 335854 366968 335860
rect 366824 335708 366876 335714
rect 366824 335650 366876 335656
rect 366088 335640 366140 335646
rect 366088 335582 366140 335588
rect 367020 7274 367048 336602
rect 367848 336530 367876 338014
rect 367836 336524 367888 336530
rect 367836 336466 367888 336472
rect 367468 336320 367520 336326
rect 367468 336262 367520 336268
rect 367008 7268 367060 7274
rect 367008 7210 367060 7216
rect 367480 6914 367508 336262
rect 368124 334490 368152 338014
rect 368216 338014 368368 338042
rect 368736 338014 368980 338042
rect 369104 338014 369348 338042
rect 369472 338014 369716 338042
rect 368112 334484 368164 334490
rect 368112 334426 368164 334432
rect 368216 7410 368244 338014
rect 368952 336734 368980 338014
rect 368296 336728 368348 336734
rect 368296 336670 368348 336676
rect 368940 336728 368992 336734
rect 368940 336670 368992 336676
rect 368204 7404 368256 7410
rect 368204 7346 368256 7352
rect 368308 7342 368336 336670
rect 369320 336462 369348 338014
rect 369308 336456 369360 336462
rect 369308 336398 369360 336404
rect 369688 7478 369716 338014
rect 369780 338014 369840 338042
rect 370208 338014 370452 338042
rect 370576 338014 370820 338042
rect 370944 338014 371188 338042
rect 371312 338014 371556 338042
rect 371680 338014 371924 338042
rect 372048 338014 372292 338042
rect 369780 336818 369808 338014
rect 369780 336790 369900 336818
rect 369872 336734 369900 336790
rect 369768 336728 369820 336734
rect 369768 336670 369820 336676
rect 369860 336728 369912 336734
rect 369860 336670 369912 336676
rect 369676 7472 369728 7478
rect 369676 7414 369728 7420
rect 368296 7336 368348 7342
rect 368296 7278 368348 7284
rect 367480 6886 368244 6914
rect 367008 5568 367060 5574
rect 367008 5510 367060 5516
rect 365812 3256 365864 3262
rect 365812 3198 365864 3204
rect 365628 2916 365680 2922
rect 365628 2858 365680 2864
rect 365824 480 365852 3198
rect 367020 480 367048 5510
rect 368216 480 368244 6886
rect 369400 3324 369452 3330
rect 369400 3266 369452 3272
rect 369412 480 369440 3266
rect 369780 2990 369808 336670
rect 370424 335986 370452 338014
rect 370504 336388 370556 336394
rect 370504 336330 370556 336336
rect 370412 335980 370464 335986
rect 370412 335922 370464 335928
rect 370516 6186 370544 336330
rect 370792 335354 370820 338014
rect 370792 335326 371096 335354
rect 370596 8968 370648 8974
rect 370596 8910 370648 8916
rect 370504 6180 370556 6186
rect 370504 6122 370556 6128
rect 369768 2984 369820 2990
rect 369768 2926 369820 2932
rect 370608 480 370636 8910
rect 371068 7546 371096 335326
rect 371056 7540 371108 7546
rect 371056 7482 371108 7488
rect 371160 3058 371188 338014
rect 371528 334558 371556 338014
rect 371792 336252 371844 336258
rect 371792 336194 371844 336200
rect 371804 335354 371832 336194
rect 371896 335850 371924 338014
rect 372264 336666 372292 338014
rect 372402 337770 372430 338028
rect 372784 338014 373028 338042
rect 373152 338014 373396 338042
rect 373520 338014 373764 338042
rect 372402 337742 372476 337770
rect 372252 336660 372304 336666
rect 372252 336602 372304 336608
rect 371884 335844 371936 335850
rect 371884 335786 371936 335792
rect 372344 335844 372396 335850
rect 372344 335786 372396 335792
rect 371804 335326 371924 335354
rect 371516 334552 371568 334558
rect 371516 334494 371568 334500
rect 371896 6254 371924 335326
rect 372356 8294 372384 335786
rect 372448 8974 372476 337742
rect 373000 335918 373028 338014
rect 373368 336598 373396 338014
rect 373356 336592 373408 336598
rect 373356 336534 373408 336540
rect 372988 335912 373040 335918
rect 372988 335854 373040 335860
rect 373736 335306 373764 338014
rect 373828 338014 373888 338042
rect 374256 338014 374500 338042
rect 374624 338014 374868 338042
rect 374992 338014 375236 338042
rect 373724 335300 373776 335306
rect 373724 335242 373776 335248
rect 373828 333878 373856 338014
rect 373908 336592 373960 336598
rect 373908 336534 373960 336540
rect 373816 333872 373868 333878
rect 373816 333814 373868 333820
rect 372436 8968 372488 8974
rect 372436 8910 372488 8916
rect 372344 8288 372396 8294
rect 372344 8230 372396 8236
rect 371884 6248 371936 6254
rect 371884 6190 371936 6196
rect 372896 4072 372948 4078
rect 372896 4014 372948 4020
rect 371700 3392 371752 3398
rect 371700 3334 371752 3340
rect 371148 3052 371200 3058
rect 371148 2994 371200 3000
rect 371712 480 371740 3334
rect 372908 480 372936 4014
rect 373920 3126 373948 336534
rect 374472 336258 374500 338014
rect 374460 336252 374512 336258
rect 374460 336194 374512 336200
rect 374644 335912 374696 335918
rect 374644 335854 374696 335860
rect 374656 333946 374684 335854
rect 374644 333940 374696 333946
rect 374644 333882 374696 333888
rect 374840 325694 374868 338014
rect 375208 332450 375236 338014
rect 375300 338014 375360 338042
rect 375728 338014 375972 338042
rect 376096 338014 376248 338042
rect 376464 338014 376616 338042
rect 376832 338014 377076 338042
rect 377200 338014 377444 338042
rect 377568 338014 377812 338042
rect 375196 332444 375248 332450
rect 375196 332386 375248 332392
rect 374840 325666 375236 325694
rect 375208 5710 375236 325666
rect 375196 5704 375248 5710
rect 375196 5646 375248 5652
rect 375300 4978 375328 338014
rect 375944 336598 375972 338014
rect 375932 336592 375984 336598
rect 375932 336534 375984 336540
rect 375472 336184 375524 336190
rect 375472 336126 375524 336132
rect 375484 16574 375512 336126
rect 376220 332382 376248 338014
rect 376588 336394 376616 338014
rect 377048 336598 377076 338014
rect 376668 336592 376720 336598
rect 376668 336534 376720 336540
rect 377036 336592 377088 336598
rect 377036 336534 377088 336540
rect 376576 336388 376628 336394
rect 376576 336330 376628 336336
rect 376208 332376 376260 332382
rect 376208 332318 376260 332324
rect 375484 16546 376524 16574
rect 375208 4950 375328 4978
rect 374092 4480 374144 4486
rect 374092 4422 374144 4428
rect 373908 3120 373960 3126
rect 373908 3062 373960 3068
rect 374104 480 374132 4422
rect 375208 3194 375236 4950
rect 375288 4140 375340 4146
rect 375288 4082 375340 4088
rect 375196 3188 375248 3194
rect 375196 3130 375248 3136
rect 375300 480 375328 4082
rect 376496 480 376524 16546
rect 376680 5778 376708 336534
rect 377416 333810 377444 338014
rect 377404 333804 377456 333810
rect 377404 333746 377456 333752
rect 376668 5772 376720 5778
rect 376668 5714 376720 5720
rect 377680 4548 377732 4554
rect 377680 4490 377732 4496
rect 377692 480 377720 4490
rect 377784 3262 377812 338014
rect 377922 337770 377950 338028
rect 378304 338014 378548 338042
rect 378672 338014 378916 338042
rect 379040 338014 379192 338042
rect 379316 338014 379468 338042
rect 379684 338014 379928 338042
rect 380052 338014 380296 338042
rect 380420 338014 380664 338042
rect 377922 337742 377996 337770
rect 377864 336592 377916 336598
rect 377864 336534 377916 336540
rect 377876 5846 377904 336534
rect 377968 5914 377996 337742
rect 378520 332314 378548 338014
rect 378888 336122 378916 338014
rect 378876 336116 378928 336122
rect 378876 336058 378928 336064
rect 378508 332308 378560 332314
rect 378508 332250 378560 332256
rect 379164 325694 379192 338014
rect 379440 332246 379468 338014
rect 379900 336530 379928 338014
rect 380268 336598 380296 338014
rect 380636 336682 380664 338014
rect 380774 337770 380802 338028
rect 381156 338014 381400 338042
rect 381524 338014 381768 338042
rect 381892 338014 382044 338042
rect 380774 337742 380848 337770
rect 380820 336818 380848 337742
rect 380820 336790 381032 336818
rect 380636 336654 380940 336682
rect 380256 336592 380308 336598
rect 380256 336534 380308 336540
rect 380716 336592 380768 336598
rect 380716 336534 380768 336540
rect 379888 336524 379940 336530
rect 379888 336466 379940 336472
rect 379428 332240 379480 332246
rect 379428 332182 379480 332188
rect 379164 325666 379468 325694
rect 378876 6248 378928 6254
rect 378876 6190 378928 6196
rect 377956 5908 378008 5914
rect 377956 5850 378008 5856
rect 377864 5840 377916 5846
rect 377864 5782 377916 5788
rect 377772 3256 377824 3262
rect 377772 3198 377824 3204
rect 378888 480 378916 6190
rect 379440 5982 379468 325666
rect 380728 6050 380756 336534
rect 380808 336524 380860 336530
rect 380808 336466 380860 336472
rect 380716 6044 380768 6050
rect 380716 5986 380768 5992
rect 379428 5976 379480 5982
rect 379428 5918 379480 5924
rect 379980 4004 380032 4010
rect 379980 3946 380032 3952
rect 379992 480 380020 3946
rect 380820 3330 380848 336466
rect 380912 333742 380940 336654
rect 381004 336326 381032 336790
rect 381372 336530 381400 338014
rect 381360 336524 381412 336530
rect 381360 336466 381412 336472
rect 381740 336394 381768 338014
rect 382016 336598 382044 338014
rect 382108 338014 382260 338042
rect 382628 338014 382872 338042
rect 382996 338014 383240 338042
rect 383364 338014 383516 338042
rect 383732 338014 383976 338042
rect 384100 338014 384344 338042
rect 384468 338014 384712 338042
rect 382004 336592 382056 336598
rect 382004 336534 382056 336540
rect 381912 336524 381964 336530
rect 381912 336466 381964 336472
rect 381728 336388 381780 336394
rect 381728 336330 381780 336336
rect 380992 336320 381044 336326
rect 380992 336262 381044 336268
rect 380900 333736 380952 333742
rect 380900 333678 380952 333684
rect 381924 325694 381952 336466
rect 381924 325666 382044 325694
rect 382016 6118 382044 325666
rect 382108 6798 382136 338014
rect 382188 336592 382240 336598
rect 382188 336534 382240 336540
rect 382096 6792 382148 6798
rect 382096 6734 382148 6740
rect 382004 6112 382056 6118
rect 382004 6054 382056 6060
rect 381176 4616 381228 4622
rect 381176 4558 381228 4564
rect 380808 3324 380860 3330
rect 380808 3266 380860 3272
rect 381188 480 381216 4558
rect 382200 3398 382228 336534
rect 382464 336184 382516 336190
rect 382464 336126 382516 336132
rect 382372 10328 382424 10334
rect 382372 10270 382424 10276
rect 382188 3392 382240 3398
rect 382188 3334 382240 3340
rect 382384 480 382412 10270
rect 382476 6914 382504 336126
rect 382844 332178 382872 338014
rect 383212 336190 383240 338014
rect 383488 336258 383516 338014
rect 383948 336462 383976 338014
rect 383936 336456 383988 336462
rect 383936 336398 383988 336404
rect 383476 336252 383528 336258
rect 383476 336194 383528 336200
rect 383200 336184 383252 336190
rect 383200 336126 383252 336132
rect 382924 335368 382976 335374
rect 382924 335310 382976 335316
rect 382832 332172 382884 332178
rect 382832 332114 382884 332120
rect 382936 10334 382964 335310
rect 384316 335170 384344 338014
rect 384684 335374 384712 338014
rect 384776 338014 384836 338042
rect 385204 338014 385356 338042
rect 385572 338014 385816 338042
rect 385940 338014 386184 338042
rect 384672 335368 384724 335374
rect 384672 335310 384724 335316
rect 384304 335164 384356 335170
rect 384304 335106 384356 335112
rect 382924 10328 382976 10334
rect 382924 10270 382976 10276
rect 382476 6886 383608 6914
rect 383580 480 383608 6886
rect 384776 6662 384804 338014
rect 384856 336456 384908 336462
rect 384856 336398 384908 336404
rect 384868 6730 384896 336398
rect 385328 332110 385356 338014
rect 385788 336025 385816 338014
rect 385774 336016 385830 336025
rect 385774 335951 385830 335960
rect 385316 332104 385368 332110
rect 385316 332046 385368 332052
rect 386156 325694 386184 338014
rect 386294 337770 386322 338028
rect 386676 338014 386920 338042
rect 387044 338014 387288 338042
rect 387412 338014 387656 338042
rect 386294 337742 386368 337770
rect 386340 330818 386368 337742
rect 386892 336705 386920 338014
rect 386878 336696 386934 336705
rect 386878 336631 386934 336640
rect 387260 336462 387288 338014
rect 387248 336456 387300 336462
rect 387248 336398 387300 336404
rect 387628 333674 387656 338014
rect 387720 338014 387780 338042
rect 388148 338014 388392 338042
rect 388516 338014 388760 338042
rect 388884 338014 389036 338042
rect 389252 338014 389496 338042
rect 389620 338014 389864 338042
rect 389988 338014 390140 338042
rect 387720 336546 387748 338014
rect 387720 336518 387840 336546
rect 387708 336456 387760 336462
rect 387708 336398 387760 336404
rect 387616 333668 387668 333674
rect 387616 333610 387668 333616
rect 386328 330812 386380 330818
rect 386328 330754 386380 330760
rect 386156 325666 386368 325694
rect 384856 6724 384908 6730
rect 384856 6666 384908 6672
rect 384764 6656 384816 6662
rect 384764 6598 384816 6604
rect 386340 6594 386368 325666
rect 386328 6588 386380 6594
rect 386328 6530 386380 6536
rect 387720 6526 387748 336398
rect 387812 336161 387840 336518
rect 388364 336462 388392 338014
rect 388352 336456 388404 336462
rect 388352 336398 388404 336404
rect 387798 336152 387854 336161
rect 387798 336087 387854 336096
rect 388444 336048 388496 336054
rect 388444 335990 388496 335996
rect 387708 6520 387760 6526
rect 387708 6462 387760 6468
rect 385960 6180 386012 6186
rect 385960 6122 386012 6128
rect 384764 4684 384816 4690
rect 384764 4626 384816 4632
rect 384776 480 384804 4626
rect 385972 480 386000 6122
rect 388260 4752 388312 4758
rect 388260 4694 388312 4700
rect 387156 3936 387208 3942
rect 387156 3878 387208 3884
rect 387168 480 387196 3878
rect 388272 480 388300 4694
rect 388456 4214 388484 335990
rect 388732 332042 388760 338014
rect 389008 335374 389036 338014
rect 389468 336462 389496 338014
rect 389088 336456 389140 336462
rect 389088 336398 389140 336404
rect 389456 336456 389508 336462
rect 389456 336398 389508 336404
rect 388996 335368 389048 335374
rect 388996 335310 389048 335316
rect 388720 332036 388772 332042
rect 388720 331978 388772 331984
rect 389100 6458 389128 336398
rect 389836 330750 389864 338014
rect 390112 335034 390140 338014
rect 390342 337770 390370 338028
rect 390724 338014 390968 338042
rect 391092 338014 391244 338042
rect 391368 338014 391612 338042
rect 391736 338014 391888 338042
rect 392104 338014 392348 338042
rect 392472 338014 392716 338042
rect 390342 337742 390416 337770
rect 390192 336456 390244 336462
rect 390192 336398 390244 336404
rect 390100 335028 390152 335034
rect 390100 334970 390152 334976
rect 389824 330744 389876 330750
rect 389824 330686 389876 330692
rect 389456 10328 389508 10334
rect 389456 10270 389508 10276
rect 389088 6452 389140 6458
rect 389088 6394 389140 6400
rect 388444 4208 388496 4214
rect 388444 4150 388496 4156
rect 389468 480 389496 10270
rect 390204 6390 390232 336398
rect 390192 6384 390244 6390
rect 390192 6326 390244 6332
rect 390388 6322 390416 337742
rect 390940 333606 390968 338014
rect 391216 336054 391244 338014
rect 391204 336048 391256 336054
rect 391204 335990 391256 335996
rect 391584 335354 391612 338014
rect 391584 335326 391704 335354
rect 390928 333600 390980 333606
rect 390928 333542 390980 333548
rect 390376 6316 390428 6322
rect 390376 6258 390428 6264
rect 391676 6254 391704 335326
rect 391860 331974 391888 338014
rect 391938 336696 391994 336705
rect 391938 336631 391994 336640
rect 391952 335102 391980 336631
rect 391940 335096 391992 335102
rect 391940 335038 391992 335044
rect 392320 334966 392348 338014
rect 392688 336462 392716 338014
rect 392826 337770 392854 338028
rect 392964 338014 393208 338042
rect 393576 338014 393820 338042
rect 393944 338014 394188 338042
rect 394312 338014 394464 338042
rect 392826 337742 392900 337770
rect 392676 336456 392728 336462
rect 392676 336398 392728 336404
rect 392308 334960 392360 334966
rect 392308 334902 392360 334908
rect 391848 331968 391900 331974
rect 391848 331910 391900 331916
rect 392872 330682 392900 337742
rect 392860 330676 392912 330682
rect 392860 330618 392912 330624
rect 391664 6248 391716 6254
rect 391664 6190 391716 6196
rect 391848 5500 391900 5506
rect 391848 5442 391900 5448
rect 390652 3868 390704 3874
rect 390652 3810 390704 3816
rect 390664 480 390692 3810
rect 391860 480 391888 5442
rect 392964 4282 392992 338014
rect 393136 336456 393188 336462
rect 393136 336398 393188 336404
rect 393148 6186 393176 336398
rect 393228 336116 393280 336122
rect 393228 336058 393280 336064
rect 393240 335374 393268 336058
rect 393228 335368 393280 335374
rect 393228 335310 393280 335316
rect 393792 334898 393820 338014
rect 393780 334892 393832 334898
rect 393780 334834 393832 334840
rect 394160 330614 394188 338014
rect 394148 330608 394200 330614
rect 394148 330550 394200 330556
rect 393136 6180 393188 6186
rect 393136 6122 393188 6128
rect 394436 4350 394464 338014
rect 394620 338014 394680 338042
rect 395048 338014 395292 338042
rect 395416 338014 395660 338042
rect 395784 338014 395936 338042
rect 396152 338014 396396 338042
rect 396520 338014 396764 338042
rect 396888 338014 397132 338042
rect 397256 338014 397408 338042
rect 397624 338014 397868 338042
rect 397992 338014 398236 338042
rect 398360 338014 398512 338042
rect 394620 333538 394648 338014
rect 394608 333532 394660 333538
rect 394608 333474 394660 333480
rect 395264 330478 395292 338014
rect 395632 335354 395660 338014
rect 395632 335326 395844 335354
rect 395252 330472 395304 330478
rect 395252 330414 395304 330420
rect 395344 5432 395396 5438
rect 395344 5374 395396 5380
rect 394424 4344 394476 4350
rect 394424 4286 394476 4292
rect 392952 4276 393004 4282
rect 392952 4218 393004 4224
rect 393044 4208 393096 4214
rect 393044 4150 393096 4156
rect 393056 480 393084 4150
rect 394240 3800 394292 3806
rect 394240 3742 394292 3748
rect 394252 480 394280 3742
rect 395356 480 395384 5374
rect 395816 4418 395844 335326
rect 395908 333470 395936 338014
rect 395896 333464 395948 333470
rect 395896 333406 395948 333412
rect 396368 331906 396396 338014
rect 396356 331900 396408 331906
rect 396356 331842 396408 331848
rect 396736 325694 396764 338014
rect 397104 334762 397132 338014
rect 397092 334756 397144 334762
rect 397092 334698 397144 334704
rect 397380 329186 397408 338014
rect 397840 335374 397868 338014
rect 397828 335368 397880 335374
rect 397828 335310 397880 335316
rect 398208 334830 398236 338014
rect 398196 334824 398248 334830
rect 398196 334766 398248 334772
rect 398484 334694 398512 338014
rect 398668 338014 398728 338042
rect 399096 338014 399340 338042
rect 399464 338014 399708 338042
rect 398564 335368 398616 335374
rect 398564 335310 398616 335316
rect 398472 334688 398524 334694
rect 398472 334630 398524 334636
rect 397368 329180 397420 329186
rect 397368 329122 397420 329128
rect 396736 325666 397132 325694
rect 396540 9036 396592 9042
rect 396540 8978 396592 8984
rect 395804 4412 395856 4418
rect 395804 4354 395856 4360
rect 396552 480 396580 8978
rect 397104 4486 397132 325666
rect 398576 4554 398604 335310
rect 398668 4622 398696 338014
rect 399312 333198 399340 338014
rect 399300 333192 399352 333198
rect 399300 333134 399352 333140
rect 399680 330886 399708 338014
rect 399818 337770 399846 338028
rect 400140 338014 400200 338042
rect 400568 338014 400812 338042
rect 400936 338014 401180 338042
rect 401304 338014 401548 338042
rect 401672 338014 401916 338042
rect 402040 338014 402284 338042
rect 402408 338014 402560 338042
rect 399818 337742 399892 337770
rect 399668 330880 399720 330886
rect 399668 330822 399720 330828
rect 398932 5296 398984 5302
rect 398932 5238 398984 5244
rect 398656 4616 398708 4622
rect 398656 4558 398708 4564
rect 398564 4548 398616 4554
rect 398564 4490 398616 4496
rect 397092 4480 397144 4486
rect 397092 4422 397144 4428
rect 397736 3732 397788 3738
rect 397736 3674 397788 3680
rect 397748 480 397776 3674
rect 398944 480 398972 5238
rect 399864 4690 399892 337742
rect 400140 333402 400168 338014
rect 400128 333396 400180 333402
rect 400128 333338 400180 333344
rect 400784 329118 400812 338014
rect 401152 335354 401180 338014
rect 401152 335326 401364 335354
rect 400772 329112 400824 329118
rect 400772 329054 400824 329060
rect 400128 5364 400180 5370
rect 400128 5306 400180 5312
rect 399852 4684 399904 4690
rect 399852 4626 399904 4632
rect 400140 480 400168 5306
rect 401336 4758 401364 335326
rect 401520 333266 401548 338014
rect 401508 333260 401560 333266
rect 401508 333202 401560 333208
rect 401888 330546 401916 338014
rect 402256 335374 402284 338014
rect 402244 335368 402296 335374
rect 402244 335310 402296 335316
rect 402532 334626 402560 338014
rect 402624 338014 402776 338042
rect 403144 338014 403296 338042
rect 403420 338014 403664 338042
rect 403788 338014 404032 338042
rect 402520 334620 402572 334626
rect 402520 334562 402572 334568
rect 401876 330540 401928 330546
rect 401876 330482 401928 330488
rect 402520 5228 402572 5234
rect 402520 5170 402572 5176
rect 401324 4752 401376 4758
rect 401324 4694 401376 4700
rect 401324 3664 401376 3670
rect 401324 3606 401376 3612
rect 401336 480 401364 3606
rect 402532 480 402560 5170
rect 402624 4078 402652 338014
rect 402704 335368 402756 335374
rect 402704 335310 402756 335316
rect 402716 5506 402744 335310
rect 402796 330540 402848 330546
rect 402796 330482 402848 330488
rect 402704 5500 402756 5506
rect 402704 5442 402756 5448
rect 402808 4146 402836 330482
rect 403268 330478 403296 338014
rect 403256 330472 403308 330478
rect 403256 330414 403308 330420
rect 403636 325694 403664 338014
rect 404004 335374 404032 338014
rect 404096 338014 404156 338042
rect 404524 338014 404768 338042
rect 404892 338014 405136 338042
rect 403992 335368 404044 335374
rect 403992 335310 404044 335316
rect 403636 325666 404032 325694
rect 404004 8226 404032 325666
rect 403992 8220 404044 8226
rect 403992 8162 404044 8168
rect 404096 5370 404124 338014
rect 404268 335368 404320 335374
rect 404268 335310 404320 335316
rect 404176 330472 404228 330478
rect 404176 330414 404228 330420
rect 404188 5438 404216 330414
rect 404176 5432 404228 5438
rect 404176 5374 404228 5380
rect 404084 5364 404136 5370
rect 404084 5306 404136 5312
rect 403624 5160 403676 5166
rect 403624 5102 403676 5108
rect 402796 4140 402848 4146
rect 402796 4082 402848 4088
rect 402612 4072 402664 4078
rect 402612 4014 402664 4020
rect 403636 480 403664 5102
rect 404280 4010 404308 335310
rect 404740 330478 404768 338014
rect 404728 330472 404780 330478
rect 404728 330414 404780 330420
rect 405108 330410 405136 338014
rect 405200 338014 405260 338042
rect 405384 338014 405628 338042
rect 405996 338014 406240 338042
rect 406364 338014 406608 338042
rect 405200 335374 405228 338014
rect 405188 335368 405240 335374
rect 405188 335310 405240 335316
rect 405096 330404 405148 330410
rect 405096 330346 405148 330352
rect 405384 8090 405412 338014
rect 405556 335368 405608 335374
rect 405556 335310 405608 335316
rect 405464 330472 405516 330478
rect 405464 330414 405516 330420
rect 405476 8158 405504 330414
rect 405464 8152 405516 8158
rect 405464 8094 405516 8100
rect 405372 8084 405424 8090
rect 405372 8026 405424 8032
rect 405568 5302 405596 335310
rect 406212 330478 406240 338014
rect 406580 335374 406608 338014
rect 406718 337770 406746 338028
rect 407040 338014 407100 338042
rect 407468 338014 407712 338042
rect 407836 338014 408080 338042
rect 408204 338014 408448 338042
rect 408572 338014 408816 338042
rect 408940 338014 409184 338042
rect 409308 338014 409552 338042
rect 406718 337742 406792 337770
rect 406568 335368 406620 335374
rect 406568 335310 406620 335316
rect 406200 330472 406252 330478
rect 406200 330414 406252 330420
rect 405648 330404 405700 330410
rect 405648 330346 405700 330352
rect 405556 5296 405608 5302
rect 405556 5238 405608 5244
rect 404268 4004 404320 4010
rect 404268 3946 404320 3952
rect 405660 3942 405688 330346
rect 406764 8022 406792 337742
rect 406844 335368 406896 335374
rect 406844 335310 406896 335316
rect 406752 8016 406804 8022
rect 406752 7958 406804 7964
rect 406856 5234 406884 335310
rect 406936 330472 406988 330478
rect 406936 330414 406988 330420
rect 406844 5228 406896 5234
rect 406844 5170 406896 5176
rect 406016 5092 406068 5098
rect 406016 5034 406068 5040
rect 405648 3936 405700 3942
rect 405648 3878 405700 3884
rect 404820 3596 404872 3602
rect 404820 3538 404872 3544
rect 404832 480 404860 3538
rect 406028 480 406056 5034
rect 406948 3874 406976 330414
rect 406936 3868 406988 3874
rect 406936 3810 406988 3816
rect 407040 3806 407068 338014
rect 407684 335374 407712 338014
rect 407672 335368 407724 335374
rect 408052 335354 408080 338014
rect 408316 335368 408368 335374
rect 408052 335326 408264 335354
rect 407672 335310 407724 335316
rect 408236 7954 408264 335326
rect 408316 335310 408368 335316
rect 408224 7948 408276 7954
rect 408224 7890 408276 7896
rect 408328 5166 408356 335310
rect 408316 5160 408368 5166
rect 408316 5102 408368 5108
rect 407212 5024 407264 5030
rect 407212 4966 407264 4972
rect 407028 3800 407080 3806
rect 407028 3742 407080 3748
rect 407224 480 407252 4966
rect 408420 3738 408448 338014
rect 408788 330478 408816 338014
rect 408776 330472 408828 330478
rect 408776 330414 408828 330420
rect 409156 325694 409184 338014
rect 409524 335374 409552 338014
rect 409616 338014 409676 338042
rect 410044 338014 410288 338042
rect 410412 338014 410656 338042
rect 409512 335368 409564 335374
rect 409512 335310 409564 335316
rect 409156 325666 409552 325694
rect 409524 7886 409552 325666
rect 409512 7880 409564 7886
rect 409512 7822 409564 7828
rect 409616 5098 409644 338014
rect 409788 335368 409840 335374
rect 409788 335310 409840 335316
rect 409696 330472 409748 330478
rect 409696 330414 409748 330420
rect 409708 5098 409736 330414
rect 409604 5092 409656 5098
rect 409604 5034 409656 5040
rect 409696 5092 409748 5098
rect 409696 5034 409748 5040
rect 409604 4956 409656 4962
rect 409604 4898 409656 4904
rect 408408 3732 408460 3738
rect 408408 3674 408460 3680
rect 408408 3528 408460 3534
rect 408408 3470 408460 3476
rect 408420 480 408448 3470
rect 409616 480 409644 4898
rect 409800 3670 409828 335310
rect 410260 330478 410288 338014
rect 410248 330472 410300 330478
rect 410248 330414 410300 330420
rect 410628 330410 410656 338014
rect 410720 338014 410780 338042
rect 410904 338014 411148 338042
rect 411516 338014 411760 338042
rect 411884 338014 412128 338042
rect 410720 335374 410748 338014
rect 410708 335368 410760 335374
rect 410708 335310 410760 335316
rect 410616 330404 410668 330410
rect 410616 330346 410668 330352
rect 410904 7750 410932 338014
rect 411076 335368 411128 335374
rect 411076 335310 411128 335316
rect 410984 330472 411036 330478
rect 410984 330414 411036 330420
rect 410996 7818 411024 330414
rect 410984 7812 411036 7818
rect 410984 7754 411036 7760
rect 410892 7744 410944 7750
rect 410892 7686 410944 7692
rect 411088 4962 411116 335310
rect 411732 330478 411760 338014
rect 412100 335374 412128 338014
rect 412238 337770 412266 338028
rect 412468 338014 412620 338042
rect 412988 338014 413232 338042
rect 413356 338014 413600 338042
rect 413724 338014 413968 338042
rect 414092 338014 414336 338042
rect 414460 338014 414704 338042
rect 412238 337742 412312 337770
rect 412088 335368 412140 335374
rect 412088 335310 412140 335316
rect 411720 330472 411772 330478
rect 411720 330414 411772 330420
rect 411168 330404 411220 330410
rect 411168 330346 411220 330352
rect 411076 4956 411128 4962
rect 411076 4898 411128 4904
rect 410800 4888 410852 4894
rect 410800 4830 410852 4836
rect 409788 3664 409840 3670
rect 409788 3606 409840 3612
rect 410812 480 410840 4830
rect 411180 3602 411208 330346
rect 412284 7682 412312 337742
rect 412364 335368 412416 335374
rect 412364 335310 412416 335316
rect 412272 7676 412324 7682
rect 412272 7618 412324 7624
rect 412376 4894 412404 335310
rect 412364 4888 412416 4894
rect 412364 4830 412416 4836
rect 411168 3596 411220 3602
rect 411168 3538 411220 3544
rect 412468 3466 412496 338014
rect 413204 335646 413232 338014
rect 413192 335640 413244 335646
rect 413192 335582 413244 335588
rect 413572 335354 413600 338014
rect 413836 335640 413888 335646
rect 413836 335582 413888 335588
rect 413572 335326 413784 335354
rect 412548 330472 412600 330478
rect 412548 330414 412600 330420
rect 412560 3534 412588 330414
rect 413756 7614 413784 335326
rect 413744 7608 413796 7614
rect 413744 7550 413796 7556
rect 413848 4826 413876 335582
rect 413100 4820 413152 4826
rect 413100 4762 413152 4768
rect 413836 4820 413888 4826
rect 413836 4762 413888 4768
rect 412548 3528 412600 3534
rect 412548 3470 412600 3476
rect 411904 3460 411956 3466
rect 411904 3402 411956 3408
rect 412456 3460 412508 3466
rect 412456 3402 412508 3408
rect 411916 480 411944 3402
rect 413112 480 413140 4762
rect 413940 3777 413968 338014
rect 414308 330478 414336 338014
rect 414676 335578 414704 338014
rect 414814 337770 414842 338028
rect 414814 337742 414888 337770
rect 414860 335646 414888 337742
rect 414848 335640 414900 335646
rect 414848 335582 414900 335588
rect 414664 335572 414716 335578
rect 414664 335514 414716 335520
rect 414296 330472 414348 330478
rect 414296 330414 414348 330420
rect 414952 20670 414980 457286
rect 416056 353258 416084 458798
rect 429844 458720 429896 458726
rect 429844 458662 429896 458668
rect 428556 458448 428608 458454
rect 428556 458390 428608 458396
rect 418804 457360 418856 457366
rect 418804 457302 418856 457308
rect 417424 457020 417476 457026
rect 417424 456962 417476 456968
rect 416044 353252 416096 353258
rect 416044 353194 416096 353200
rect 415124 335640 415176 335646
rect 415124 335582 415176 335588
rect 414940 20664 414992 20670
rect 414940 20606 414992 20612
rect 414296 7064 414348 7070
rect 414296 7006 414348 7012
rect 413926 3768 413982 3777
rect 413926 3703 413982 3712
rect 414308 480 414336 7006
rect 415136 3369 415164 335582
rect 415308 335572 415360 335578
rect 415308 335514 415360 335520
rect 415216 330472 415268 330478
rect 415216 330414 415268 330420
rect 415228 3505 415256 330414
rect 415320 3641 415348 335514
rect 416780 335504 416832 335510
rect 416780 335446 416832 335452
rect 416792 4162 416820 335446
rect 417436 167006 417464 456962
rect 418816 405686 418844 457302
rect 425704 457292 425756 457298
rect 425704 457234 425756 457240
rect 421656 457156 421708 457162
rect 421656 457098 421708 457104
rect 418804 405680 418856 405686
rect 418804 405622 418856 405628
rect 421564 335640 421616 335646
rect 421564 335582 421616 335588
rect 418160 335436 418212 335442
rect 418160 335378 418212 335384
rect 417424 167000 417476 167006
rect 417424 166942 417476 166948
rect 418172 16574 418200 335378
rect 418804 335368 418856 335374
rect 418804 335310 418856 335316
rect 418172 16546 418752 16574
rect 417884 7132 417936 7138
rect 417884 7074 417936 7080
rect 416700 4134 416820 4162
rect 415306 3632 415362 3641
rect 415306 3567 415362 3576
rect 415214 3496 415270 3505
rect 415214 3431 415270 3440
rect 415122 3360 415178 3369
rect 415122 3295 415178 3304
rect 415492 2848 415544 2854
rect 415492 2790 415544 2796
rect 415504 480 415532 2790
rect 416700 480 416728 4134
rect 417896 480 417924 7074
rect 418724 3482 418752 16546
rect 418816 4214 418844 335310
rect 421576 8362 421604 335582
rect 421668 273222 421696 457098
rect 425716 379506 425744 457234
rect 425704 379500 425756 379506
rect 425704 379442 425756 379448
rect 425704 335844 425756 335850
rect 425704 335786 425756 335792
rect 425060 335708 425112 335714
rect 425060 335650 425112 335656
rect 421656 273216 421708 273222
rect 421656 273158 421708 273164
rect 421564 8356 421616 8362
rect 421564 8298 421616 8304
rect 423772 8356 423824 8362
rect 423772 8298 423824 8304
rect 421380 7200 421432 7206
rect 421380 7142 421432 7148
rect 418804 4208 418856 4214
rect 418804 4150 418856 4156
rect 420184 4208 420236 4214
rect 420184 4150 420236 4156
rect 418724 3454 419028 3482
rect 419000 480 419028 3454
rect 420196 480 420224 4150
rect 421392 480 421420 7142
rect 422576 2916 422628 2922
rect 422576 2858 422628 2864
rect 422588 480 422616 2858
rect 423784 480 423812 8298
rect 424968 7268 425020 7274
rect 424968 7210 425020 7216
rect 424980 480 425008 7210
rect 425072 6914 425100 335650
rect 425716 7342 425744 335786
rect 428464 335776 428516 335782
rect 428464 335718 428516 335724
rect 428476 8362 428504 335718
rect 428568 325650 428596 458390
rect 429856 431934 429884 458662
rect 432604 458584 432656 458590
rect 432604 458526 432656 458532
rect 431224 456952 431276 456958
rect 431224 456894 431276 456900
rect 429844 431928 429896 431934
rect 429844 431870 429896 431876
rect 429200 335912 429252 335918
rect 429200 335854 429252 335860
rect 428556 325644 428608 325650
rect 428556 325586 428608 325592
rect 429212 16574 429240 335854
rect 430580 334484 430632 334490
rect 430580 334426 430632 334432
rect 430592 16574 430620 334426
rect 431236 20670 431264 456894
rect 432616 365702 432644 458526
rect 432604 365696 432656 365702
rect 432604 365638 432656 365644
rect 436100 336728 436152 336734
rect 436100 336670 436152 336676
rect 432602 336152 432658 336161
rect 432602 336087 432658 336096
rect 431224 20664 431276 20670
rect 431224 20606 431276 20612
rect 429212 16546 429700 16574
rect 430592 16546 430896 16574
rect 428464 8356 428516 8362
rect 428464 8298 428516 8304
rect 425704 7336 425756 7342
rect 425704 7278 425756 7284
rect 427268 7336 427320 7342
rect 427268 7278 427320 7284
rect 425072 6886 425744 6914
rect 425716 3482 425744 6886
rect 425716 3454 426204 3482
rect 426176 480 426204 3454
rect 427280 480 427308 7278
rect 428464 7268 428516 7274
rect 428464 7210 428516 7216
rect 428476 480 428504 7210
rect 429672 480 429700 16546
rect 430868 480 430896 16546
rect 432616 9042 432644 336087
rect 435364 335980 435416 335986
rect 435364 335922 435416 335928
rect 432604 9036 432656 9042
rect 432604 8978 432656 8984
rect 434444 8356 434496 8362
rect 434444 8298 434496 8304
rect 432052 7404 432104 7410
rect 432052 7346 432104 7352
rect 432064 480 432092 7346
rect 433248 2984 433300 2990
rect 433248 2926 433300 2932
rect 433260 480 433288 2926
rect 434456 480 434484 8298
rect 435376 7546 435404 335922
rect 436112 16574 436140 336670
rect 443000 336660 443052 336666
rect 443000 336602 443052 336608
rect 440332 334552 440384 334558
rect 440332 334494 440384 334500
rect 436112 16546 436784 16574
rect 435364 7540 435416 7546
rect 435364 7482 435416 7488
rect 435548 7336 435600 7342
rect 435548 7278 435600 7284
rect 435560 480 435588 7278
rect 436756 480 436784 16546
rect 437940 7540 437992 7546
rect 437940 7482 437992 7488
rect 437952 480 437980 7482
rect 439136 7404 439188 7410
rect 439136 7346 439188 7352
rect 439148 480 439176 7346
rect 440344 3058 440372 334494
rect 443012 16574 443040 336602
rect 449900 336592 449952 336598
rect 449900 336534 449952 336540
rect 448520 335300 448572 335306
rect 448520 335242 448572 335248
rect 445760 333940 445812 333946
rect 445760 333882 445812 333888
rect 445772 16574 445800 333882
rect 443012 16546 443868 16574
rect 445772 16546 446260 16574
rect 442632 8288 442684 8294
rect 442632 8230 442684 8236
rect 440240 3052 440292 3058
rect 440240 2994 440292 3000
rect 440332 3052 440384 3058
rect 440332 2994 440384 3000
rect 441528 3052 441580 3058
rect 441528 2994 441580 3000
rect 440252 1578 440280 2994
rect 440252 1550 440372 1578
rect 440344 480 440372 1550
rect 441540 480 441568 2994
rect 442644 480 442672 8230
rect 443840 480 443868 16546
rect 445024 8968 445076 8974
rect 445024 8910 445076 8916
rect 445036 480 445064 8910
rect 446232 480 446260 16546
rect 448532 6914 448560 335242
rect 448612 333872 448664 333878
rect 448612 333814 448664 333820
rect 448624 11762 448652 333814
rect 449912 16574 449940 336534
rect 456800 336524 456852 336530
rect 456800 336466 456852 336472
rect 452660 332444 452712 332450
rect 452660 332386 452712 332392
rect 452672 16574 452700 332386
rect 449912 16546 450952 16574
rect 452672 16546 453344 16574
rect 448612 11756 448664 11762
rect 448612 11698 448664 11704
rect 449808 11756 449860 11762
rect 449808 11698 449860 11704
rect 448532 6886 448652 6914
rect 447416 3120 447468 3126
rect 447416 3062 447468 3068
rect 447428 480 447456 3062
rect 448624 480 448652 6886
rect 449820 480 449848 11698
rect 450924 480 450952 16546
rect 452108 5704 452160 5710
rect 452108 5646 452160 5652
rect 452120 480 452148 5646
rect 453316 480 453344 16546
rect 455696 5772 455748 5778
rect 455696 5714 455748 5720
rect 454500 3188 454552 3194
rect 454500 3130 454552 3136
rect 454512 480 454540 3130
rect 455708 480 455736 5714
rect 456812 1426 456840 336466
rect 465080 336456 465132 336462
rect 465080 336398 465132 336404
rect 459560 333804 459612 333810
rect 459560 333746 459612 333752
rect 456892 332376 456944 332382
rect 456892 332318 456944 332324
rect 456800 1420 456852 1426
rect 456800 1362 456852 1368
rect 456904 480 456932 332318
rect 459572 16574 459600 333746
rect 463700 332308 463752 332314
rect 463700 332250 463752 332256
rect 463712 16574 463740 332250
rect 465092 16574 465120 336398
rect 468484 336388 468536 336394
rect 468484 336330 468536 336336
rect 466460 332240 466512 332246
rect 466460 332182 466512 332188
rect 466472 16574 466500 332182
rect 459572 16546 460428 16574
rect 463712 16546 464016 16574
rect 465092 16546 465212 16574
rect 466472 16546 467512 16574
rect 459192 5840 459244 5846
rect 459192 5782 459244 5788
rect 458088 1420 458140 1426
rect 458088 1362 458140 1368
rect 458100 480 458128 1362
rect 459204 480 459232 5782
rect 460400 480 460428 16546
rect 462780 5908 462832 5914
rect 462780 5850 462832 5856
rect 461584 3256 461636 3262
rect 461584 3198 461636 3204
rect 461596 480 461624 3198
rect 462792 480 462820 5850
rect 463988 480 464016 16546
rect 465184 480 465212 16546
rect 466276 5976 466328 5982
rect 466276 5918 466328 5924
rect 466288 480 466316 5918
rect 467484 480 467512 16546
rect 468496 5982 468524 336330
rect 471980 336320 472032 336326
rect 471980 336262 472032 336268
rect 470600 333736 470652 333742
rect 470600 333678 470652 333684
rect 470612 16574 470640 333678
rect 471992 16574 472020 336262
rect 475384 336252 475436 336258
rect 475384 336194 475436 336200
rect 470612 16546 471100 16574
rect 471992 16546 472296 16574
rect 469864 6044 469916 6050
rect 469864 5986 469916 5992
rect 468484 5976 468536 5982
rect 468484 5918 468536 5924
rect 468668 3324 468720 3330
rect 468668 3266 468720 3272
rect 468680 480 468708 3266
rect 469876 480 469904 5986
rect 471072 480 471100 16546
rect 472268 480 472296 16546
rect 473452 6112 473504 6118
rect 473452 6054 473504 6060
rect 473464 480 473492 6054
rect 474556 5976 474608 5982
rect 474556 5918 474608 5924
rect 474568 480 474596 5918
rect 475396 5574 475424 336194
rect 478880 336184 478932 336190
rect 478880 336126 478932 336132
rect 477500 332172 477552 332178
rect 477500 332114 477552 332120
rect 477512 16574 477540 332114
rect 478892 16574 478920 336126
rect 497464 336116 497516 336122
rect 497464 336058 497516 336064
rect 486422 336016 486478 336025
rect 486422 335951 486478 335960
rect 483020 335232 483072 335238
rect 483020 335174 483072 335180
rect 481640 335164 481692 335170
rect 481640 335106 481692 335112
rect 477512 16546 478184 16574
rect 478892 16546 479380 16574
rect 476948 6792 477000 6798
rect 476948 6734 477000 6740
rect 475384 5568 475436 5574
rect 475384 5510 475436 5516
rect 475752 3392 475804 3398
rect 475752 3334 475804 3340
rect 475764 480 475792 3334
rect 476960 480 476988 6734
rect 478156 480 478184 16546
rect 479352 480 479380 16546
rect 480536 5568 480588 5574
rect 480536 5510 480588 5516
rect 480548 480 480576 5510
rect 481652 3398 481680 335106
rect 483032 16574 483060 335174
rect 485780 332104 485832 332110
rect 485780 332046 485832 332052
rect 485044 330880 485096 330886
rect 485044 330822 485096 330828
rect 483032 16546 484072 16574
rect 481732 6724 481784 6730
rect 481732 6666 481784 6672
rect 481640 3392 481692 3398
rect 481640 3334 481692 3340
rect 481744 480 481772 6666
rect 482836 3392 482888 3398
rect 482836 3334 482888 3340
rect 482848 480 482876 3334
rect 484044 480 484072 16546
rect 485056 3330 485084 330822
rect 485792 6914 485820 332046
rect 486436 16574 486464 335951
rect 490012 335096 490064 335102
rect 490012 335038 490064 335044
rect 489184 330812 489236 330818
rect 489184 330754 489236 330760
rect 486436 16546 486556 16574
rect 485792 6886 486464 6914
rect 485228 6656 485280 6662
rect 485228 6598 485280 6604
rect 485044 3324 485096 3330
rect 485044 3266 485096 3272
rect 485240 480 485268 6598
rect 486436 480 486464 6886
rect 486528 5574 486556 16546
rect 488816 6588 488868 6594
rect 488816 6530 488868 6536
rect 486516 5568 486568 5574
rect 486516 5510 486568 5516
rect 487620 5568 487672 5574
rect 487620 5510 487672 5516
rect 487632 480 487660 5510
rect 488828 480 488856 6530
rect 489196 3398 489224 330754
rect 490024 16574 490052 335038
rect 492680 333668 492732 333674
rect 492680 333610 492732 333616
rect 492692 16574 492720 333610
rect 496820 332036 496872 332042
rect 496820 331978 496872 331984
rect 496832 16574 496860 331978
rect 490024 16546 491156 16574
rect 492692 16546 493548 16574
rect 496832 16546 497136 16574
rect 489184 3392 489236 3398
rect 489184 3334 489236 3340
rect 489920 3392 489972 3398
rect 489920 3334 489972 3340
rect 489932 480 489960 3334
rect 491128 480 491156 16546
rect 492312 6520 492364 6526
rect 492312 6462 492364 6468
rect 492324 480 492352 6462
rect 493520 480 493548 16546
rect 494704 9036 494756 9042
rect 494704 8978 494756 8984
rect 494716 480 494744 8978
rect 495900 6452 495952 6458
rect 495900 6394 495952 6400
rect 495912 480 495940 6394
rect 497108 480 497136 16546
rect 497476 5574 497504 336058
rect 504364 336048 504416 336054
rect 504364 335990 504416 335996
rect 500960 335028 501012 335034
rect 500960 334970 501012 334976
rect 499580 330744 499632 330750
rect 499580 330686 499632 330692
rect 499592 16574 499620 330686
rect 500972 16574 501000 334970
rect 502984 333600 503036 333606
rect 502984 333542 503036 333548
rect 499592 16546 500632 16574
rect 500972 16546 501828 16574
rect 499396 6384 499448 6390
rect 499396 6326 499448 6332
rect 497464 5568 497516 5574
rect 497464 5510 497516 5516
rect 498200 5568 498252 5574
rect 498200 5510 498252 5516
rect 498212 480 498240 5510
rect 499408 480 499436 6326
rect 500604 480 500632 16546
rect 501800 480 501828 16546
rect 502892 6316 502944 6322
rect 502892 6258 502944 6264
rect 502904 3210 502932 6258
rect 502996 3330 503024 333542
rect 504376 5574 504404 335990
rect 507860 334960 507912 334966
rect 507860 334902 507912 334908
rect 506480 331968 506532 331974
rect 506480 331910 506532 331916
rect 504364 5568 504416 5574
rect 504364 5510 504416 5516
rect 505376 5568 505428 5574
rect 505376 5510 505428 5516
rect 502984 3324 503036 3330
rect 502984 3266 503036 3272
rect 504180 3324 504232 3330
rect 504180 3266 504232 3272
rect 502904 3182 503024 3210
rect 502996 480 503024 3182
rect 504192 480 504220 3266
rect 505388 480 505416 5510
rect 506492 3330 506520 331910
rect 507872 16574 507900 334902
rect 512644 334892 512696 334898
rect 512644 334834 512696 334840
rect 510620 330676 510672 330682
rect 510620 330618 510672 330624
rect 510632 16574 510660 330618
rect 507872 16546 508912 16574
rect 510632 16546 511304 16574
rect 506572 6248 506624 6254
rect 506572 6190 506624 6196
rect 506480 3324 506532 3330
rect 506480 3266 506532 3272
rect 506584 3210 506612 6190
rect 507676 3324 507728 3330
rect 507676 3266 507728 3272
rect 506492 3182 506612 3210
rect 506492 480 506520 3182
rect 507688 480 507716 3266
rect 508884 480 508912 16546
rect 510068 6180 510120 6186
rect 510068 6122 510120 6128
rect 510080 480 510108 6122
rect 511276 480 511304 16546
rect 512460 4276 512512 4282
rect 512460 4218 512512 4224
rect 512472 480 512500 4218
rect 512656 3194 512684 334834
rect 526444 334824 526496 334830
rect 526444 334766 526496 334772
rect 522304 334756 522356 334762
rect 522304 334698 522356 334704
rect 515404 333532 515456 333538
rect 515404 333474 515456 333480
rect 514760 330608 514812 330614
rect 514760 330550 514812 330556
rect 512644 3188 512696 3194
rect 512644 3130 512696 3136
rect 513564 3188 513616 3194
rect 513564 3130 513616 3136
rect 513576 480 513604 3130
rect 514772 480 514800 330550
rect 515416 3330 515444 333474
rect 520280 333464 520332 333470
rect 520280 333406 520332 333412
rect 519544 331900 519596 331906
rect 519544 331842 519596 331848
rect 517520 330540 517572 330546
rect 517520 330482 517572 330488
rect 517532 16574 517560 330482
rect 519556 16574 519584 331842
rect 520292 16574 520320 333406
rect 517532 16546 518388 16574
rect 519556 16546 519676 16574
rect 520292 16546 520780 16574
rect 515956 4344 516008 4350
rect 515956 4286 516008 4292
rect 515404 3324 515456 3330
rect 515404 3266 515456 3272
rect 515968 480 515996 4286
rect 517152 3324 517204 3330
rect 517152 3266 517204 3272
rect 517164 480 517192 3266
rect 518360 480 518388 16546
rect 519544 4412 519596 4418
rect 519544 4354 519596 4360
rect 519556 480 519584 4354
rect 519648 3330 519676 16546
rect 519636 3324 519688 3330
rect 519636 3266 519688 3272
rect 520752 480 520780 16546
rect 522316 3330 522344 334698
rect 524420 329180 524472 329186
rect 524420 329122 524472 329128
rect 524432 16574 524460 329122
rect 524432 16546 525472 16574
rect 523040 4480 523092 4486
rect 523040 4422 523092 4428
rect 521844 3324 521896 3330
rect 521844 3266 521896 3272
rect 522304 3324 522356 3330
rect 522304 3266 522356 3272
rect 521856 480 521884 3266
rect 523052 480 523080 4422
rect 524236 3324 524288 3330
rect 524236 3266 524288 3272
rect 524248 480 524276 3266
rect 525444 480 525472 16546
rect 526456 3262 526484 334766
rect 528560 334688 528612 334694
rect 528560 334630 528612 334636
rect 528572 16574 528600 334630
rect 540244 334620 540296 334626
rect 540244 334562 540296 334568
rect 530584 333396 530636 333402
rect 530584 333338 530636 333344
rect 528572 16546 529060 16574
rect 526628 4548 526680 4554
rect 526628 4490 526680 4496
rect 526444 3256 526496 3262
rect 526444 3198 526496 3204
rect 526640 480 526668 4490
rect 527824 3256 527876 3262
rect 527824 3198 527876 3204
rect 527836 480 527864 3198
rect 529032 480 529060 16546
rect 530124 4616 530176 4622
rect 530124 4558 530176 4564
rect 530136 480 530164 4558
rect 530596 3398 530624 333338
rect 533344 333328 533396 333334
rect 533344 333270 533396 333276
rect 533356 3398 533384 333270
rect 538220 333260 538272 333266
rect 538220 333202 538272 333208
rect 535460 329112 535512 329118
rect 535460 329054 535512 329060
rect 535472 16574 535500 329054
rect 538232 16574 538260 333202
rect 535472 16546 536144 16574
rect 538232 16546 538444 16574
rect 533712 4684 533764 4690
rect 533712 4626 533764 4632
rect 530584 3392 530636 3398
rect 530584 3334 530636 3340
rect 531320 3392 531372 3398
rect 531320 3334 531372 3340
rect 533344 3392 533396 3398
rect 533344 3334 533396 3340
rect 531332 480 531360 3334
rect 532516 3324 532568 3330
rect 532516 3266 532568 3272
rect 532528 480 532556 3266
rect 533724 480 533752 4626
rect 534908 3392 534960 3398
rect 534908 3334 534960 3340
rect 534920 480 534948 3334
rect 536116 480 536144 16546
rect 537208 4752 537260 4758
rect 537208 4694 537260 4700
rect 537220 480 537248 4694
rect 538416 480 538444 16546
rect 540256 3398 540284 334562
rect 562336 259418 562364 459546
rect 566476 313274 566504 459614
rect 569236 419490 569264 459682
rect 580264 458312 580316 458318
rect 580264 458254 580316 458260
rect 579802 458144 579858 458153
rect 579802 458079 579858 458088
rect 579816 456890 579844 458079
rect 579804 456884 579856 456890
rect 579804 456826 579856 456832
rect 580172 431928 580224 431934
rect 580172 431870 580224 431876
rect 580184 431633 580212 431870
rect 580170 431624 580226 431633
rect 580170 431559 580226 431568
rect 569224 419484 569276 419490
rect 569224 419426 569276 419432
rect 580172 419484 580224 419490
rect 580172 419426 580224 419432
rect 580184 418305 580212 419426
rect 580170 418296 580226 418305
rect 580170 418231 580226 418240
rect 579620 405680 579672 405686
rect 579620 405622 579672 405628
rect 579632 404977 579660 405622
rect 579618 404968 579674 404977
rect 579618 404903 579674 404912
rect 580172 379500 580224 379506
rect 580172 379442 580224 379448
rect 580184 378457 580212 379442
rect 580170 378448 580226 378457
rect 580170 378383 580226 378392
rect 580172 365696 580224 365702
rect 580172 365638 580224 365644
rect 580184 365129 580212 365638
rect 580170 365120 580226 365129
rect 580170 365055 580226 365064
rect 580172 353252 580224 353258
rect 580172 353194 580224 353200
rect 580184 351937 580212 353194
rect 580170 351928 580226 351937
rect 580170 351863 580226 351872
rect 579896 325644 579948 325650
rect 579896 325586 579948 325592
rect 579908 325281 579936 325586
rect 579894 325272 579950 325281
rect 579894 325207 579950 325216
rect 566464 313268 566516 313274
rect 566464 313210 566516 313216
rect 580172 313268 580224 313274
rect 580172 313210 580224 313216
rect 580184 312089 580212 313210
rect 580170 312080 580226 312089
rect 580170 312015 580226 312024
rect 580276 298761 580304 458254
rect 580262 298752 580318 298761
rect 580262 298687 580318 298696
rect 580172 273216 580224 273222
rect 580172 273158 580224 273164
rect 580184 272241 580212 273158
rect 580170 272232 580226 272241
rect 580170 272167 580226 272176
rect 562324 259412 562376 259418
rect 562324 259354 562376 259360
rect 580172 259412 580224 259418
rect 580172 259354 580224 259360
rect 580184 258913 580212 259354
rect 580170 258904 580226 258913
rect 580170 258839 580226 258848
rect 580172 167000 580224 167006
rect 580172 166942 580224 166948
rect 580184 165889 580212 166942
rect 580170 165880 580226 165889
rect 580170 165815 580226 165824
rect 579988 20664 580040 20670
rect 579988 20606 580040 20612
rect 580000 19825 580028 20606
rect 579986 19816 580042 19825
rect 579986 19751 580042 19760
rect 545488 8220 545540 8226
rect 545488 8162 545540 8168
rect 540796 5500 540848 5506
rect 540796 5442 540848 5448
rect 539600 3392 539652 3398
rect 539600 3334 539652 3340
rect 540244 3392 540296 3398
rect 540244 3334 540296 3340
rect 539612 480 539640 3334
rect 540808 480 540836 5442
rect 544384 5432 544436 5438
rect 544384 5374 544436 5380
rect 543188 4072 543240 4078
rect 543188 4014 543240 4020
rect 541992 3392 542044 3398
rect 541992 3334 542044 3340
rect 542004 480 542032 3334
rect 543200 480 543228 4014
rect 544396 480 544424 5374
rect 545500 480 545528 8162
rect 549076 8152 549128 8158
rect 549076 8094 549128 8100
rect 547880 5364 547932 5370
rect 547880 5306 547932 5312
rect 546684 4004 546736 4010
rect 546684 3946 546736 3952
rect 546696 480 546724 3946
rect 547892 480 547920 5306
rect 549088 480 549116 8094
rect 552664 8084 552716 8090
rect 552664 8026 552716 8032
rect 551468 5296 551520 5302
rect 551468 5238 551520 5244
rect 550272 3936 550324 3942
rect 550272 3878 550324 3884
rect 550284 480 550312 3878
rect 551480 480 551508 5238
rect 552676 480 552704 8026
rect 556160 8016 556212 8022
rect 556160 7958 556212 7964
rect 554964 5228 555016 5234
rect 554964 5170 555016 5176
rect 553768 3868 553820 3874
rect 553768 3810 553820 3816
rect 553780 480 553808 3810
rect 554976 480 555004 5170
rect 556172 480 556200 7958
rect 559748 7948 559800 7954
rect 559748 7890 559800 7896
rect 558552 5160 558604 5166
rect 558552 5102 558604 5108
rect 557356 3800 557408 3806
rect 557356 3742 557408 3748
rect 557368 480 557396 3742
rect 558564 480 558592 5102
rect 559760 480 559788 7890
rect 56t 412